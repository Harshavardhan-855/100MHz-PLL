magic
tech sky130A
timestamp 1709124411
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
use inverter  x1
timestamp 1709123519
transform 1 0 202 0 1 -754
box -202 154 395 781
use inverter  x2
timestamp 1709123519
transform 1 0 799 0 1 -754
box -202 154 395 781
use inverteraaa  x3aaa
timestamp 1709123519
transform 1 0 1396 0 1 -754
box -202 154 395 781
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 inp
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 out
port 3 nsew
<< end >>
