magic
tech sky130A
magscale 1 2
timestamp 1713428059
<< error_p >>
rect -29 161 29 167
rect -29 127 -17 161
rect -29 121 29 127
rect -29 -127 29 -121
rect -29 -161 -17 -127
rect -29 -167 29 -161
<< nwell >>
rect -211 -299 211 299
<< pmos >>
rect -15 -80 15 80
<< pdiff >>
rect -73 51 -15 80
rect -73 17 -61 51
rect -27 17 -15 51
rect -73 -17 -15 17
rect -73 -51 -61 -17
rect -27 -51 -15 -17
rect -73 -80 -15 -51
rect 15 51 73 80
rect 15 17 27 51
rect 61 17 73 51
rect 15 -17 73 17
rect 15 -51 27 -17
rect 61 -51 73 -17
rect 15 -80 73 -51
<< pdiffc >>
rect -61 17 -27 51
rect -61 -51 -27 -17
rect 27 17 61 51
rect 27 -51 61 -17
<< nsubdiff >>
rect -175 229 -51 263
rect -17 229 17 263
rect 51 229 175 263
rect -175 153 -141 229
rect -175 85 -141 119
rect 141 153 175 229
rect 141 85 175 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -119 -141 -85
rect -175 -229 -141 -153
rect 141 -119 175 -85
rect 141 -229 175 -153
rect -175 -263 -51 -229
rect -17 -263 17 -229
rect 51 -263 175 -229
<< nsubdiffcont >>
rect -51 229 -17 263
rect 17 229 51 263
rect -175 119 -141 153
rect 141 119 175 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -153 -141 -119
rect 141 -153 175 -119
rect -51 -263 -17 -229
rect 17 -263 51 -229
<< poly >>
rect -33 161 33 177
rect -33 127 -17 161
rect 17 127 33 161
rect -33 111 33 127
rect -15 80 15 111
rect -15 -111 15 -80
rect -33 -127 33 -111
rect -33 -161 -17 -127
rect 17 -161 33 -127
rect -33 -177 33 -161
<< polycont >>
rect -17 127 17 161
rect -17 -161 17 -127
<< locali >>
rect -175 229 -51 263
rect -17 229 17 263
rect 51 229 175 263
rect -175 153 -141 229
rect -33 127 -17 161
rect 17 127 33 161
rect 141 153 175 229
rect -175 85 -141 119
rect 141 85 175 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -61 53 -27 84
rect -61 -17 -27 17
rect -61 -84 -27 -53
rect 27 53 61 84
rect 27 -17 61 17
rect 27 -84 61 -53
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -119 -141 -85
rect 141 -119 175 -85
rect -175 -229 -141 -153
rect -33 -161 -17 -127
rect 17 -161 33 -127
rect 141 -229 175 -153
rect -175 -263 -51 -229
rect -17 -263 17 -229
rect 51 -263 175 -229
<< viali >>
rect -17 127 17 161
rect -61 51 -27 53
rect -61 19 -27 51
rect -61 -51 -27 -19
rect -61 -53 -27 -51
rect 27 51 61 53
rect 27 19 61 51
rect 27 -51 61 -19
rect 27 -53 61 -51
rect -17 -161 17 -127
<< metal1 >>
rect -29 161 29 167
rect -29 127 -17 161
rect 17 127 29 161
rect -29 121 29 127
rect -67 53 -21 80
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -80 -21 -53
rect 21 53 67 80
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -80 67 -53
rect -29 -127 29 -121
rect -29 -161 -17 -127
rect 17 -161 29 -127
rect -29 -167 29 -161
<< properties >>
string FIXED_BBOX -158 -246 158 246
<< end >>
