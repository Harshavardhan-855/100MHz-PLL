magic
tech sky130A
magscale 1 2
timestamp 1713431446
<< nwell >>
rect 3896 5068 3964 5234
rect 3924 4948 4008 4990
rect 3838 4746 4008 4948
rect 3838 4728 4006 4746
rect 4068 3726 4100 3828
rect 3476 2734 3492 2738
rect 3476 2728 3798 2734
<< pwell >>
rect 1600 4380 1642 4384
rect 990 4210 1142 4368
rect 1600 4152 1646 4380
rect 1986 4152 2158 4182
rect 1600 4108 2158 4152
rect 1602 4106 2158 4108
rect 998 3362 1150 3520
rect 1600 3302 1678 3522
rect 1600 3240 2134 3302
rect 1600 3238 1678 3240
rect 990 2536 1142 2694
rect 1588 2390 1668 2680
<< locali >>
rect 1030 5350 2062 5442
rect 2164 5434 4264 5444
rect 2164 5378 4274 5434
rect 4080 5326 4274 5378
rect 4080 5276 4084 5326
rect 4002 5214 4084 5276
rect 1358 5114 1504 5162
rect 2358 5124 2504 5172
rect 2846 5112 2992 5160
rect 3266 5114 3412 5162
rect 3686 5120 3832 5168
rect 4000 5150 4084 5214
rect 4126 4498 4272 5148
rect 1026 4316 1142 4368
rect 1026 4272 1150 4316
rect 1026 4268 1148 4272
rect 1026 4210 1142 4268
rect 4116 3938 4272 4498
rect 4116 3928 4268 3938
rect 4126 3652 4268 3928
rect 1022 3464 1150 3520
rect 1022 3420 1154 3464
rect 1022 3362 1150 3420
rect 1718 3194 1828 3534
rect 4116 3082 4268 3652
rect 4120 3080 4268 3082
rect 4120 2810 4266 3080
rect 3742 2712 4266 2810
rect 1018 2616 1142 2682
rect 3434 2664 3476 2668
rect 3434 2630 3438 2664
rect 3472 2630 3476 2664
rect 3434 2626 3476 2630
rect 3742 2628 3778 2712
rect 1018 2572 1152 2616
rect 1018 2524 1142 2572
rect 3110 2440 3234 2480
rect 3432 2382 3480 2570
rect 3900 2382 4078 2422
rect 3430 2296 4078 2382
<< viali >>
rect 838 5146 1030 5442
rect 4084 5148 4276 5326
rect 850 4108 1026 4568
rect 846 3222 1022 3682
rect 854 2478 1018 2850
rect 3438 2630 3472 2664
rect 3898 2422 4080 2600
<< metal1 >>
rect 1158 5480 1358 5680
rect 832 5442 1036 5454
rect 832 5146 838 5442
rect 1030 5146 1036 5442
rect 832 5134 1036 5146
rect 1188 5310 1314 5480
rect 2160 5324 3896 5330
rect 1188 5258 1916 5310
rect 2152 5262 3896 5324
rect 4072 5326 4288 5332
rect 838 4594 1030 5134
rect 1188 5024 1314 5258
rect 2152 5168 2210 5262
rect 3920 5234 3996 5238
rect 1930 5110 2308 5168
rect 3074 5108 3160 5228
rect 3506 5108 3564 5226
rect 3896 5108 3996 5234
rect 4072 5148 4084 5326
rect 4276 5148 4288 5326
rect 4072 5142 4288 5148
rect 4084 5130 4284 5142
rect 3082 5106 3170 5108
rect 3506 5106 3574 5108
rect 3044 5080 3170 5106
rect 1188 4972 1918 5024
rect 834 4568 1034 4594
rect 834 4108 850 4568
rect 1026 4108 1034 4568
rect 834 3682 1034 4108
rect 834 3222 846 3682
rect 1022 3222 1034 3682
rect 834 2850 1034 3222
rect 834 2478 854 2850
rect 1018 2526 1034 2850
rect 1018 2478 1040 2526
rect 834 2340 1040 2478
rect 1188 2443 1314 4972
rect 2298 4970 2364 5020
rect 2984 4970 3050 5020
rect 3082 4700 3170 5080
rect 3462 5078 3574 5106
rect 3890 5080 4006 5108
rect 3406 4968 3472 5018
rect 3506 4922 3574 5078
rect 3896 5068 4006 5080
rect 3828 4970 3894 5020
rect 3922 4990 4006 5068
rect 3922 4924 4008 4990
rect 3426 4770 3436 4922
rect 3594 4770 3604 4922
rect 3830 4742 3840 4924
rect 4000 4742 4010 4924
rect 3136 4698 3170 4700
rect 1880 4468 1934 4672
rect 3128 4664 3162 4698
rect 2908 4580 2956 4610
rect 4026 4604 4076 4670
rect 1600 4380 1642 4384
rect 1600 4152 1646 4380
rect 1860 4358 1870 4468
rect 2106 4358 2116 4468
rect 2762 4400 2956 4580
rect 2762 4398 4088 4400
rect 1880 4182 1934 4358
rect 2762 4326 4092 4398
rect 2762 4244 2956 4326
rect 2908 4242 2956 4244
rect 3006 4182 3056 4248
rect 1986 4164 2158 4182
rect 1968 4152 2158 4164
rect 1600 4150 1720 4152
rect 1756 4150 2158 4152
rect 1600 4108 2158 4150
rect 1602 4106 2158 4108
rect 1882 3666 1936 3824
rect 3378 3812 3388 3888
rect 3706 3812 3716 3888
rect 4026 3828 4092 4326
rect 4026 3824 4100 3828
rect 2912 3750 2958 3764
rect 1874 3576 1884 3666
rect 2072 3576 2082 3666
rect 1600 3414 1678 3522
rect 1576 3378 1690 3414
rect 1600 3302 1678 3378
rect 1882 3330 1936 3576
rect 2678 3556 2958 3750
rect 4012 3738 4100 3824
rect 4012 3576 4028 3738
rect 4018 3572 4028 3576
rect 4090 3572 4100 3738
rect 2678 3468 3504 3556
rect 2678 3462 3288 3468
rect 2678 3394 2958 3462
rect 2912 3392 2958 3394
rect 3010 3332 3060 3398
rect 1728 3302 1764 3314
rect 1984 3302 2014 3322
rect 1600 3240 2134 3302
rect 1600 3238 1678 3240
rect 1726 3236 2014 3240
rect 1880 3082 1890 3202
rect 2184 3082 2194 3202
rect 3278 3188 3288 3462
rect 3502 3320 3512 3468
rect 3502 3314 4024 3320
rect 3502 3198 4114 3314
rect 3502 3188 3512 3198
rect 1886 2978 1944 3082
rect 1882 2854 1944 2978
rect 3312 2962 3322 3052
rect 3982 2962 3992 3052
rect 2910 2914 2956 2916
rect 2768 2860 2956 2914
rect 4026 2910 4114 3198
rect 1588 2458 1668 2680
rect 1882 2486 1934 2854
rect 2768 2610 2778 2860
rect 2942 2836 2956 2860
rect 2942 2790 3486 2836
rect 2942 2772 2956 2790
rect 2942 2694 2954 2772
rect 2942 2610 2956 2694
rect 3436 2674 3486 2790
rect 3422 2664 3488 2674
rect 3422 2630 3438 2664
rect 3472 2630 3488 2664
rect 3422 2620 3488 2630
rect 2768 2548 2956 2610
rect 3886 2600 4092 2606
rect 3008 2486 3058 2552
rect 1588 2388 2252 2458
rect 3886 2422 3898 2600
rect 4080 2422 4092 2600
rect 3886 2416 4092 2422
rect 3892 2404 4092 2416
rect 840 2326 1040 2340
<< via1 >>
rect 3436 4770 3594 4922
rect 3840 4742 4000 4924
rect 1870 4358 2106 4468
rect 3388 3812 3706 3888
rect 1884 3576 2072 3666
rect 4028 3572 4090 3738
rect 1890 3082 2184 3202
rect 3288 3188 3502 3468
rect 3322 2962 3982 3052
rect 2778 2610 2942 2860
<< metal2 >>
rect 3436 4922 3594 4932
rect 3436 4760 3594 4770
rect 3838 4924 4006 4948
rect 1870 4468 2106 4478
rect 2106 4358 2372 4466
rect 1870 4356 2372 4358
rect 1870 4348 2106 4356
rect 1884 3666 2072 3676
rect 1884 3566 2072 3576
rect 1890 3202 2184 3212
rect 1890 3072 2184 3082
rect 2258 2768 2370 4356
rect 3436 3898 3592 4760
rect 3838 4742 3840 4924
rect 4000 4742 4006 4924
rect 3838 4728 4006 4742
rect 3388 3888 3706 3898
rect 3388 3802 3706 3812
rect 3288 3468 3502 3478
rect 3838 3476 3982 4728
rect 4028 3738 4090 3748
rect 4028 3562 4090 3572
rect 3702 3470 3982 3476
rect 3288 3178 3502 3188
rect 3700 3062 3982 3470
rect 3322 3052 3982 3062
rect 3322 2952 3982 2962
rect 2778 2860 2942 2870
rect 2258 2698 2778 2768
rect 2258 2694 2370 2698
rect 2778 2600 2942 2610
<< via2 >>
rect 1884 3576 2072 3666
rect 1890 3082 2184 3202
rect 4028 3572 4090 3738
rect 3288 3188 3502 3468
<< metal3 >>
rect 4018 3738 4100 3743
rect 1874 3668 2082 3671
rect 4018 3668 4028 3738
rect 1874 3666 4028 3668
rect 1874 3576 1884 3666
rect 2072 3576 4028 3666
rect 1874 3574 4028 3576
rect 1874 3571 2082 3574
rect 4018 3572 4028 3574
rect 4090 3572 4100 3738
rect 4018 3567 4100 3572
rect 3278 3468 3512 3473
rect 3278 3232 3288 3468
rect 1900 3207 3288 3232
rect 1880 3202 3288 3207
rect 1880 3082 1890 3202
rect 2184 3188 3288 3202
rect 3502 3188 3512 3468
rect 2184 3183 3512 3188
rect 2184 3098 3498 3183
rect 2184 3082 2194 3098
rect 1880 3077 2194 3082
use sky130_fd_pr__nfet_01v8_MMRDEV  M1
timestamp 1713428059
transform -1 0 1718 0 -1 5140
box -386 -280 386 280
use sky130_fd_pr__pfet_01v8_XYUFBL  M2
timestamp 1713428059
transform 1 0 2331 0 1 5147
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XYUFBL  M3
timestamp 1713428059
transform 1 0 3439 0 1 5145
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  M4
timestamp 1713428059
transform 0 1 2981 -1 0 3789
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  M5
timestamp 1713428059
transform 1 0 1366 0 1 3444
box -386 -280 386 280
use sky130_fd_pr__nfet_01v8_BBNS5X  M6
timestamp 1713428059
transform 0 1 2472 -1 0 3365
box -201 -700 201 700
use sky130_fd_pr__pfet_01v8_XYUFBL  M7
timestamp 1713428059
transform 1 0 3861 0 1 5147
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  M8
timestamp 1713428059
transform 0 1 2981 -1 0 2943
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  M9
timestamp 1713428059
transform -1 0 1364 0 1 2596
box -386 -280 386 280
use sky130_fd_pr__nfet_01v8_BBNS5X  M10
timestamp 1713428059
transform 0 1 2470 1 0 2519
box -201 -700 201 700
use sky130_fd_pr__pfet_01v8_XYUFBL  M11
timestamp 1713428059
transform 1 0 3017 0 1 5147
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  M12
timestamp 1713428059
transform 0 1 2979 -1 0 4637
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  M13
timestamp 1713428059
transform 1 0 1362 0 1 4292
box -386 -280 386 280
use sky130_fd_pr__nfet_01v8_BBNS5X  M14
timestamp 1713428059
transform 0 1 2468 -1 0 4215
box -201 -700 201 700
use sky130_fd_sc_hd__inv_2  x1
timestamp 1713428059
transform 0 1 3216 -1 0 2692
box -38 -48 314 592
<< labels >>
flabel metal1 s 3892 2404 4092 2604 0 FreeSans 320 0 0 0 out
port 4 nsew
flabel metal1 s 4084 5130 4284 5330 0 FreeSans 320 180 0 0 vdd
port 1 nsew
flabel metal1 s 840 2326 1040 2526 0 FreeSans 320 0 0 0 vss
port 2 nsew
flabel metal1 s 1158 5480 1358 5680 0 FreeSans 320 0 0 0 vctrl
port 3 nsew
<< end >>
