magic
tech sky130A
magscale 1 2
timestamp 1713418706
<< nwell >>
rect 3704 374 3908 384
rect 3672 328 3908 374
rect 3704 44 3908 328
rect 2376 -702 2832 -372
rect 3426 -696 3632 -370
rect 3674 -1434 3858 -1116
<< pwell >>
rect 3656 -150 3894 -14
rect 2360 -934 2862 -762
rect 3368 -892 3610 -760
rect 3610 -1674 3834 -1480
<< psubdiff >>
rect 3694 -148 3718 -18
rect 3870 -148 3894 -18
rect 3434 -882 3458 -786
rect 3584 -882 3608 -786
rect 3704 -1502 3834 -1478
rect 3704 -1700 3834 -1676
<< nsubdiff >>
rect 3708 311 3796 338
rect 3708 217 3737 311
rect 3771 217 3796 311
rect 3708 198 3796 217
rect 3710 192 3796 198
rect 3498 -471 3586 -444
rect 3498 -565 3527 -471
rect 3561 -565 3586 -471
rect 3498 -584 3586 -565
rect 3500 -590 3586 -584
rect 3690 -1179 3778 -1152
rect 3690 -1273 3719 -1179
rect 3753 -1273 3778 -1179
rect 3690 -1292 3778 -1273
rect 3692 -1298 3778 -1292
<< psubdiffcont >>
rect 3718 -148 3870 -18
rect 3458 -882 3584 -786
rect 3704 -1676 3834 -1502
<< nsubdiffcont >>
rect 3737 217 3771 311
rect 3527 -565 3561 -471
rect 3719 -1273 3753 -1179
<< locali >>
rect 3658 312 3772 346
rect 1750 256 1814 312
rect 3737 311 3771 312
rect 3737 196 3771 217
rect 890 104 1560 106
rect 942 -16 1560 104
rect 3702 -48 3718 -18
rect 3870 -48 3886 -18
rect 3884 -146 3886 -48
rect 3702 -148 3718 -146
rect 3870 -148 3886 -146
rect 3294 -430 3558 -388
rect 3484 -436 3558 -430
rect 3484 -470 3562 -436
rect 3527 -471 3561 -470
rect 3527 -586 3561 -565
rect 1852 -780 1982 -662
rect 2282 -752 2648 -702
rect 2816 -744 3012 -692
rect 3338 -738 4078 -626
rect 2816 -746 2836 -744
rect 2964 -746 3012 -744
rect 1704 -1226 1766 -1168
rect 3548 -1172 3756 -1134
rect 3674 -1178 3754 -1172
rect 3719 -1179 3753 -1178
rect 3719 -1294 3753 -1273
rect 878 -1502 1470 -1374
rect 3704 -1502 3834 -1486
<< viali >>
rect 752 -18 942 104
rect 3312 8 3376 122
rect 3698 -146 3718 -48
rect 3718 -146 3870 -48
rect 3870 -146 3884 -48
rect 1706 -790 1852 -656
rect 2648 -754 2816 -690
rect 3142 -740 3210 -678
rect 4078 -750 4288 -572
rect 3438 -786 3606 -776
rect 3438 -882 3458 -786
rect 3458 -882 3584 -786
rect 3584 -882 3606 -786
rect 3438 -886 3606 -882
rect 712 -1508 878 -1372
rect 3266 -1494 3324 -1366
rect 3700 -1676 3704 -1522
rect 3704 -1676 3834 -1522
rect 3834 -1676 3836 -1522
rect 3700 -1704 3836 -1676
<< metal1 >>
rect 1132 378 1374 608
rect 1132 280 1534 378
rect 696 110 896 154
rect 696 104 954 110
rect 696 -18 752 104
rect 942 -18 954 104
rect 696 -24 954 -18
rect 696 -46 896 -24
rect 1132 -340 1374 280
rect 3306 132 3382 134
rect 4054 132 4254 162
rect 3306 122 4254 132
rect 3306 8 3312 122
rect 3376 8 4254 122
rect 3306 4 4254 8
rect 3306 -4 3382 4
rect 2421 -94 2431 -28
rect 2523 -94 2533 -28
rect 4054 -38 4254 4
rect 3658 -48 3966 -42
rect 3658 -146 3698 -48
rect 3884 -146 3966 -48
rect 3658 -166 3966 -146
rect 3644 -264 3968 -166
rect 1122 -488 1132 -340
rect 1360 -374 1374 -340
rect 1908 -374 1918 -372
rect 1360 -474 1918 -374
rect 2116 -470 2126 -372
rect 2330 -468 2890 -360
rect 1360 -488 1374 -474
rect 1132 -1106 1374 -488
rect 1694 -656 1864 -650
rect 1694 -790 1706 -656
rect 1852 -790 1864 -656
rect 3130 -678 3222 -672
rect 2636 -690 2828 -684
rect 3130 -688 3142 -678
rect 2636 -698 2648 -690
rect 2634 -754 2648 -698
rect 2816 -754 2828 -690
rect 2636 -760 2828 -754
rect 3122 -756 3132 -688
rect 3210 -740 3222 -678
rect 3200 -746 3222 -740
rect 3200 -756 3210 -746
rect 3702 -752 3968 -264
rect 4076 -566 4236 -38
rect 3610 -758 3968 -752
rect 4066 -572 4300 -566
rect 4066 -750 4078 -572
rect 4288 -750 4300 -572
rect 4066 -756 4300 -750
rect 1694 -796 1864 -790
rect 3394 -776 3968 -758
rect 3394 -886 3438 -776
rect 3606 -886 3968 -776
rect 2933 -908 3007 -906
rect 3394 -908 3968 -886
rect 2354 -1016 3968 -908
rect 1132 -1200 1474 -1106
rect 1132 -1208 1374 -1200
rect 3610 -1202 3640 -1102
rect 656 -1366 856 -1330
rect 3260 -1366 3330 -1354
rect 656 -1372 890 -1366
rect 656 -1508 712 -1372
rect 878 -1508 890 -1372
rect 3260 -1494 3266 -1366
rect 3324 -1368 3666 -1366
rect 3324 -1492 3562 -1368
rect 3654 -1492 3666 -1368
rect 3324 -1494 3330 -1492
rect 3260 -1506 3330 -1494
rect 656 -1514 890 -1508
rect 3702 -1510 3968 -1016
rect 4124 -1336 4324 -1308
rect 4094 -1352 4324 -1336
rect 4014 -1502 4024 -1352
rect 4098 -1502 4324 -1352
rect 4124 -1508 4324 -1502
rect 656 -1530 856 -1514
rect 2502 -1566 2512 -1512
rect 2602 -1566 2612 -1512
rect 3694 -1522 3968 -1510
rect 3694 -1648 3700 -1522
rect 3628 -1704 3700 -1648
rect 3836 -1704 3968 -1522
rect 3628 -1746 3968 -1704
rect 3702 -1968 3968 -1746
<< via1 >>
rect 2431 -94 2523 -28
rect 1132 -488 1360 -340
rect 1918 -470 2116 -372
rect 1706 -790 1852 -656
rect 3132 -740 3142 -688
rect 3142 -740 3200 -688
rect 3132 -756 3200 -740
rect 3562 -1492 3654 -1368
rect 4024 -1502 4098 -1352
rect 2512 -1566 2602 -1512
<< metal2 >>
rect 2431 -28 2523 -18
rect 2429 -94 2431 -28
rect 2429 -104 2523 -94
rect 1706 -264 1848 -262
rect 2429 -264 2521 -104
rect 1132 -340 1360 -330
rect 1132 -498 1360 -488
rect 1706 -332 2522 -264
rect 1706 -614 1848 -332
rect 1918 -372 2116 -362
rect 1918 -480 2116 -470
rect 1704 -646 1848 -614
rect 1704 -656 1852 -646
rect 1704 -790 1706 -656
rect 3132 -688 3200 -678
rect 1704 -800 1852 -790
rect 3126 -756 3132 -690
rect 3200 -756 3202 -690
rect 1704 -1034 1840 -800
rect 1702 -1100 2602 -1034
rect 3126 -1046 3202 -756
rect 3126 -1092 3648 -1046
rect 2514 -1502 2602 -1100
rect 3568 -1358 3648 -1092
rect 4024 -1352 4098 -1342
rect 3562 -1362 3654 -1358
rect 3562 -1368 4024 -1362
rect 3654 -1492 4024 -1368
rect 3562 -1496 4024 -1492
rect 3562 -1502 3654 -1496
rect 2512 -1512 2602 -1502
rect 4024 -1512 4098 -1502
rect 2512 -1576 2602 -1566
use sky130_fd_sc_hd__dfrbp_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 1478 0 1 -216
box -38 -48 2246 592
use sky130_fd_sc_hd__and2_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform -1 0 3406 0 1 -956
box -38 -48 590 592
use sky130_fd_sc_hd__dfrbp_2  x3
timestamp 1712078602
transform 1 0 1432 0 1 -1698
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_4  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform -1 0 2372 0 1 -966
box -38 -48 498 592
<< labels >>
flabel metal1 3734 -1940 3934 -1740 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 656 -1530 856 -1330 0 FreeSans 256 0 0 0 B
port 5 nsew
flabel metal1 4124 -1508 4324 -1308 0 FreeSans 256 0 0 0 QB
port 4 nsew
flabel metal1 4054 -38 4254 162 0 FreeSans 256 0 0 0 QA
port 3 nsew
flabel metal1 696 -46 896 154 0 FreeSans 256 0 0 0 A
port 2 nsew
flabel metal1 1160 394 1360 594 0 FreeSans 256 0 0 0 VDD
port 1 nsew
<< end >>
