magic
tech sky130A
magscale 1 2
timestamp 1708514189
<< error_s >>
rect 2401 -264 2561 -262
rect 2429 -292 2533 -290
rect 2429 -346 2943 -332
rect 2429 -348 2533 -346
rect 2401 -374 2943 -360
rect 2401 -376 2561 -374
rect 2837 -691 2845 -632
rect 2871 -657 2879 -607
rect 2837 -818 2845 -745
rect 2871 -852 2879 -779
rect 2421 -1012 2619 -1004
rect 2421 -1016 2933 -1012
rect 2449 -1040 2591 -1032
rect 2449 -1044 2933 -1040
rect 2449 -1084 3007 -1078
rect 2449 -1088 2591 -1084
rect 2421 -1112 3035 -1106
rect 2421 -1116 2619 -1112
rect 2423 -1474 2617 -1462
rect 2451 -1502 2589 -1490
<< locali >>
rect 1750 256 1814 312
rect 890 104 1560 106
rect 942 -16 1560 104
rect 1704 -1226 1766 -1168
rect 878 -1502 1470 -1374
<< viali >>
rect 752 -18 942 104
rect 3312 8 3376 122
rect 2777 -818 2845 -632
rect 712 -1508 878 -1372
rect 3266 -1494 3324 -1366
<< metal1 >>
rect 1132 378 1374 608
rect 1132 280 1534 378
rect 696 110 896 154
rect 696 104 954 110
rect 696 -18 752 104
rect 942 -18 954 104
rect 696 -24 954 -18
rect 696 -46 896 -24
rect 1132 -340 1374 280
rect 3306 132 3382 134
rect 4054 132 4254 162
rect 3306 122 4254 132
rect 3306 8 3312 122
rect 3376 8 4254 122
rect 3306 4 4254 8
rect 3306 -4 3382 4
rect 2421 -94 2431 -28
rect 2523 -94 2533 -28
rect 4054 -38 4254 4
rect 3644 -264 3968 -166
rect 1122 -488 1132 -340
rect 1360 -488 1374 -340
rect 2429 -348 2439 -290
rect 2523 -296 2533 -290
rect 2523 -300 3003 -296
rect 2523 -346 3007 -300
rect 2523 -348 2533 -346
rect 2943 -360 3007 -346
rect 1908 -470 1918 -372
rect 2116 -470 2126 -372
rect 2330 -468 3007 -360
rect 1132 -1106 1374 -488
rect 2771 -632 2851 -620
rect 2771 -698 2777 -632
rect 2266 -754 2777 -698
rect 2771 -818 2777 -754
rect 2845 -660 2851 -632
rect 2943 -660 3007 -468
rect 2845 -790 3007 -660
rect 2845 -818 2851 -790
rect 2771 -830 2851 -818
rect 2933 -908 3007 -790
rect 3702 -908 3968 -264
rect 2354 -1016 3968 -908
rect 2449 -1088 2459 -1032
rect 2581 -1040 2591 -1032
rect 2933 -1040 3007 -1016
rect 2581 -1084 3007 -1040
rect 2581 -1088 2591 -1084
rect 1132 -1200 1474 -1106
rect 1132 -1208 1374 -1200
rect 3610 -1202 3640 -1102
rect 656 -1366 856 -1330
rect 3260 -1366 3330 -1354
rect 656 -1372 890 -1366
rect 656 -1508 712 -1372
rect 878 -1508 890 -1372
rect 656 -1514 890 -1508
rect 656 -1530 856 -1514
rect 2451 -1546 2461 -1490
rect 2579 -1546 2589 -1490
rect 3260 -1494 3266 -1366
rect 3324 -1368 3666 -1366
rect 3324 -1492 3562 -1368
rect 3654 -1492 3666 -1368
rect 3324 -1494 3330 -1492
rect 3260 -1506 3330 -1494
rect 3702 -1648 3968 -1016
rect 4124 -1336 4324 -1308
rect 4094 -1352 4324 -1336
rect 4014 -1502 4024 -1352
rect 4098 -1502 4324 -1352
rect 4124 -1508 4324 -1502
rect 3628 -1746 3968 -1648
rect 3702 -1968 3968 -1746
<< via1 >>
rect 2431 -94 2523 -28
rect 1132 -488 1360 -340
rect 2439 -348 2523 -290
rect 1918 -470 2116 -372
rect 2459 -1088 2581 -1032
rect 2461 -1546 2579 -1490
rect 3562 -1492 3654 -1368
rect 4024 -1502 4098 -1352
<< metal2 >>
rect 2431 -28 2523 -18
rect 2429 -94 2431 -28
rect 2429 -104 2523 -94
rect 2429 -280 2521 -104
rect 2429 -290 2523 -280
rect 1132 -340 1360 -330
rect 2429 -334 2439 -290
rect 2439 -358 2523 -348
rect 1918 -372 2116 -362
rect 1360 -470 1918 -374
rect 1360 -474 2116 -470
rect 1918 -480 2116 -474
rect 1132 -498 1360 -488
rect 2459 -1032 2581 -1022
rect 2459 -1098 2581 -1088
rect 2465 -1480 2579 -1098
rect 4024 -1352 4098 -1342
rect 2461 -1490 2579 -1480
rect 3562 -1362 3654 -1358
rect 3562 -1368 4024 -1362
rect 3654 -1492 4024 -1368
rect 3562 -1496 4024 -1492
rect 3562 -1502 3654 -1496
rect 4024 -1512 4098 -1502
rect 2461 -1556 2579 -1546
use sky130_fd_sc_hd__dfrbp_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform 1 0 1478 0 1 -216
box -38 -48 2246 592
use sky130_fd_sc_hd__and2_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform -1 0 3406 0 1 -956
box -38 -48 590 592
use sky130_fd_sc_hd__dfrbp_2  x3
timestamp 1705271942
transform 1 0 1432 0 1 -1698
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_4  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform -1 0 2372 0 1 -966
box -38 -48 498 592
<< labels >>
flabel metal1 1160 394 1360 594 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 3734 -1940 3934 -1740 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 696 -46 896 154 0 FreeSans 256 0 0 0 A
port 2 nsew
flabel metal1 656 -1530 856 -1330 0 FreeSans 256 0 0 0 B
port 5 nsew
flabel metal1 4054 -38 4254 162 0 FreeSans 256 0 0 0 QA
port 3 nsew
flabel metal1 4124 -1508 4324 -1308 0 FreeSans 256 0 0 0 QB
port 4 nsew
<< end >>
