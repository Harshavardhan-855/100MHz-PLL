magic
tech sky130A
magscale 1 2
timestamp 1713443771
<< pwell >>
rect 11466 -1336 11496 -1326
<< psubdiff >>
rect 11466 -1336 11496 -1326
<< locali >>
rect 3398 1966 3402 2018
rect 3592 1964 3840 2016
rect 4137 1949 4346 2009
rect -20 426 332 592
rect -20 -20 -16 426
rect 330 -20 332 426
rect 5476 -760 6004 -746
rect 5476 -808 5644 -760
rect 5474 -1336 5644 -808
rect 11466 -1336 11496 -1326
rect 5474 -1938 5916 -1336
<< viali >>
rect 3402 1942 3592 2078
rect 4346 1904 4470 2028
rect -16 -22 330 426
rect 5644 -1336 6104 -760
rect 7058 -1336 11374 -1184
rect 11500 -1850 11788 -1310
<< metal1 >>
rect 4582 2706 4856 2956
rect 504 2558 4502 2572
rect 504 2386 3748 2558
rect 4486 2386 4502 2558
rect 504 2346 4502 2386
rect 504 2318 3754 2346
rect 3000 2250 3754 2318
rect 4352 2318 4502 2346
rect 4352 2250 4362 2318
rect 3000 2248 4354 2250
rect 20 1902 266 2174
rect 4622 2154 4822 2706
rect 4904 2572 6858 2594
rect 4904 2400 4926 2572
rect 5664 2416 6858 2572
rect 9566 2436 9576 2698
rect 9828 2436 9838 2698
rect 5664 2400 6874 2416
rect 4904 2390 6874 2400
rect 4904 2376 6226 2390
rect 4904 2294 4914 2376
rect 6216 2290 6226 2294
rect 6504 2290 6874 2390
rect 3390 2078 3604 2084
rect 3390 1942 3402 2078
rect 3592 1942 3604 2078
rect 6322 2074 6874 2290
rect 4618 2034 4628 2046
rect 3390 1936 3604 1942
rect 4334 2028 4628 2034
rect 4334 1904 4346 2028
rect 4470 1904 4628 2028
rect 4334 1898 4628 1904
rect 4618 1836 4628 1898
rect 4722 2034 4732 2046
rect 4722 1898 4762 2034
rect 4722 1836 4732 1898
rect 3044 1544 3054 1802
rect 3308 1544 3318 1802
rect 3748 1704 3758 1800
rect 3998 1704 4008 1800
rect 6224 1300 6234 1792
rect 6544 1300 6554 1792
rect 4624 1266 4842 1280
rect 4622 1158 4632 1266
rect 4826 1158 4842 1266
rect -64 653 336 660
rect -67 451 336 653
rect -64 426 336 451
rect -64 -22 -16 426
rect 330 -22 336 426
rect -64 -30 336 -22
rect -22 -34 336 -30
rect 476 68 718 1061
rect 4622 1042 4842 1158
rect 3458 846 4628 1042
rect 4828 846 4842 1042
rect 3458 842 4842 846
rect 4624 840 4842 842
rect 6004 721 6230 722
rect 6295 721 6561 1069
rect 6004 495 6563 721
rect 6004 488 6230 495
rect 3046 222 6230 488
rect 476 -22 3512 68
rect 35 -1720 237 -34
rect 476 -638 718 -22
rect 476 -728 3519 -638
rect 5650 -702 5660 -260
rect 5866 -702 5876 -260
rect 476 -1338 718 -728
rect 6004 -748 6230 222
rect 6854 -632 6864 -418
rect 7066 -632 7076 -418
rect 5638 -760 6230 -748
rect 5638 -1336 5644 -760
rect 6104 -785 6230 -760
rect 9918 -785 10120 -534
rect 11398 -772 12086 -766
rect 11398 -785 11530 -772
rect 6104 -1184 11530 -785
rect 6104 -1336 7058 -1184
rect 11374 -1278 11530 -1184
rect 12078 -1278 12088 -772
rect 11374 -1310 12086 -1278
rect 11374 -1336 11500 -1310
rect 476 -1428 3519 -1338
rect 5638 -1348 6110 -1336
rect 7046 -1342 11386 -1336
rect 476 -1430 718 -1428
rect 35 -1922 3258 -1720
rect 6238 -1728 6248 -1428
rect 6718 -1728 6728 -1428
rect 10948 -1726 10958 -1418
rect 11412 -1726 11422 -1418
rect 11494 -1850 11500 -1336
rect 11788 -1326 12086 -1310
rect 11788 -1850 11794 -1326
rect 11494 -1862 11794 -1850
rect 11523 -2585 11789 -1862
<< via1 >>
rect 3748 2386 4486 2558
rect 3754 2250 4352 2346
rect 4926 2400 5664 2572
rect 9576 2436 9828 2698
rect 6226 2376 6504 2390
rect 4914 2294 6504 2376
rect 6226 2290 6504 2294
rect 4628 1836 4722 2046
rect 3054 1544 3308 1802
rect 3758 1704 3998 1800
rect 6234 1300 6544 1792
rect 4632 1158 4826 1266
rect 4628 846 4828 1042
rect 5660 -702 5866 -260
rect 6864 -632 7066 -418
rect 11530 -1278 12078 -772
rect 6248 -1728 6718 -1428
rect 10958 -1726 11412 -1418
<< metal2 >>
rect 9576 2698 9828 2708
rect 3704 2572 5710 2594
rect 3704 2558 4926 2572
rect 3704 2386 3748 2558
rect 4486 2400 4926 2558
rect 5664 2400 5710 2572
rect 9576 2426 9828 2436
rect 4486 2386 5710 2400
rect 6226 2390 6504 2400
rect 3704 2376 6226 2386
rect 3704 2370 4914 2376
rect 3738 2346 4914 2370
rect 3738 2284 3754 2346
rect 4352 2294 4914 2346
rect 4352 2290 6226 2294
rect 6504 2290 6506 2380
rect 4352 2284 6506 2290
rect 6226 2280 6504 2284
rect 3754 2240 4352 2250
rect 4628 2048 4722 2056
rect 4626 2046 4826 2048
rect 4626 1836 4628 2046
rect 4722 1836 4826 2046
rect 4628 1826 4722 1836
rect 3054 1802 3308 1812
rect 3758 1800 3998 1810
rect 3308 1704 3758 1798
rect 3308 1698 3998 1704
rect 3758 1694 3998 1698
rect 6234 1792 6544 1802
rect 3054 1534 3308 1544
rect 6234 1290 6544 1300
rect 4632 1266 4826 1276
rect 4826 1158 4832 1258
rect 4632 1052 4832 1158
rect 4628 1042 4832 1052
rect 4828 934 4832 1042
rect 4628 836 4828 846
rect 5654 -176 5966 -166
rect 5966 -418 7074 -398
rect 5966 -632 6864 -418
rect 7066 -632 7074 -418
rect 5966 -672 7074 -632
rect 5654 -722 5966 -712
rect 11530 -772 12078 -762
rect 11530 -1288 12078 -1278
rect 10958 -1418 11412 -1408
rect 6248 -1428 6718 -1418
rect 6248 -1738 6718 -1728
rect 10958 -1736 11412 -1726
<< via2 >>
rect 9576 2436 9828 2698
rect 6234 1300 6544 1792
rect 5654 -260 5966 -176
rect 5654 -702 5660 -260
rect 5660 -702 5866 -260
rect 5866 -702 5966 -260
rect 5654 -712 5966 -702
rect 11530 -1278 12078 -772
rect 6248 -1728 6718 -1428
rect 10958 -1726 11412 -1418
<< metal3 >>
rect 5654 -171 5976 3409
rect 9566 2698 9838 2703
rect 9566 2436 9576 2698
rect 9828 2436 9838 2698
rect 9566 2431 9838 2436
rect 6248 1798 6554 1800
rect 6214 1298 6224 1798
rect 6612 1298 6622 1798
rect 6224 1295 6604 1298
rect 5644 -176 5976 -171
rect 5644 -712 5654 -176
rect 5966 -712 5976 -176
rect 5644 -717 5976 -712
rect 6248 -1423 6604 1295
rect 11494 -1272 11504 -750
rect 12248 -1272 12258 -750
rect 11510 -1278 11530 -1272
rect 12078 -1278 12088 -1272
rect 11510 -1283 12088 -1278
rect 10948 -1418 11422 -1413
rect 6238 -1428 6728 -1423
rect 6238 -1728 6248 -1428
rect 6718 -1728 6728 -1428
rect 6238 -1733 6728 -1728
rect 10948 -1726 10958 -1418
rect 11412 -1726 11422 -1418
rect 10948 -1731 11422 -1726
rect 11510 -2448 12082 -1283
rect 17202 -2448 17212 -2442
rect 5464 -2454 11360 -2448
rect 5412 -2590 5422 -2454
rect 6224 -2582 11360 -2454
rect 12236 -2580 17212 -2448
rect 18218 -2580 18228 -2442
rect 12236 -2582 18194 -2580
rect 6224 -2590 6234 -2582
<< via3 >>
rect 9576 2436 9828 2698
rect 6224 1792 6612 1798
rect 6224 1300 6234 1792
rect 6234 1300 6544 1792
rect 6544 1300 6612 1792
rect 6224 1298 6612 1300
rect 11504 -772 12248 -750
rect 11504 -1272 11530 -772
rect 11530 -1272 12078 -772
rect 12078 -1272 12248 -772
rect 10958 -1726 11412 -1418
rect 5422 -2590 6224 -2454
rect 11360 -2582 12236 -2448
rect 17212 -2580 18218 -2442
<< metal4 >>
rect 9578 5532 16130 5724
rect 9578 2890 9770 5532
rect 12180 5090 12372 5532
rect 15938 5124 16130 5532
rect 9564 2698 9836 2890
rect 9564 2436 9576 2698
rect 9828 2436 9836 2698
rect 9564 2434 9836 2436
rect 9576 2420 9828 2434
rect 9576 1814 9806 2420
rect 6272 1799 10130 1814
rect 6223 1798 10130 1799
rect 6223 1298 6224 1798
rect 6612 1312 10130 1798
rect 6612 1298 6613 1312
rect 6223 1297 6613 1298
rect 11503 -750 12249 -749
rect 11503 -1272 11504 -750
rect 12248 -772 12249 -750
rect 12248 -889 12506 -772
rect 14874 -889 14996 -642
rect 19896 -889 20064 -606
rect 12248 -1130 20064 -889
rect 12248 -1147 20027 -1130
rect 12248 -1272 12506 -1147
rect 11503 -1273 12506 -1272
rect 12216 -1308 12506 -1273
rect 10957 -1418 11413 -1417
rect 10957 -1726 10958 -1418
rect 11412 -1426 11413 -1418
rect 11412 -1726 11416 -1426
rect 10957 -1727 11416 -1726
rect 10974 -2122 11416 -1727
rect 2300 -2372 15076 -2122
rect 2300 -2676 2404 -2372
rect 5421 -2454 6225 -2453
rect 5421 -2590 5422 -2454
rect 6224 -2590 6225 -2454
rect 5421 -2591 6225 -2590
rect 8632 -2666 8736 -2372
rect 11359 -2448 12237 -2447
rect 11359 -2582 11360 -2448
rect 12236 -2582 12237 -2448
rect 11359 -2583 12237 -2582
rect 14964 -2666 15068 -2372
rect 17211 -2442 18219 -2441
rect 17211 -2580 17212 -2442
rect 18218 -2580 18219 -2442
rect 17211 -2581 18219 -2580
use CHARGE_PUMP  CHARGE_PUMP_0 ~/pll/magic/cp
timestamp 1713421724
transform 1 0 4342 0 1 1012
box 280 -140 2222 1346
use divider_3N  divider_3N_0 ~/pll/magic/divider
timestamp 1713423503
transform -1 0 7450 0 1 -340
box 1588 -1636 4358 410
use pfd  pfd_0 ~/pll/magic/pfd
timestamp 1713423889
transform 1 0 -656 0 1 1968
box 656 -1746 4338 608
use sky130_fd_pr__cap_mim_m3_1_NJY377  sky130_fd_pr__cap_mim_m3_1_NJY377_0
timestamp 1713442013
transform 1 0 15094 0 1 2378
box -4892 -3040 4892 3040
use sky130_fd_pr__cap_mim_m3_1_XQ7TVA  sky130_fd_pr__cap_mim_m3_1_XQ7TVA_0
timestamp 1713432778
transform 1 0 8830 0 1 -11682
box -9378 -9120 9378 9120
use sky130_fd_pr__res_xhigh_po_1p41_K2QYT8  sky130_fd_pr__res_xhigh_po_1p41_K2QYT8_0
timestamp 1713432778
transform 0 1 8842 -1 0 -1585
box -307 -2724 307 2724
use sky130_fd_sc_hd__inv_4#0  sky130_fd_sc_hd__inv_4_0
timestamp 1712816020
transform 1 0 3756 0 1 1752
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 4216 0 1 1752
box -38 -48 130 592
use VCO_Final  VCO_Final_0 ~/pll/magic/vco
timestamp 1713431446
transform -1 0 10956 0 1 -3036
box 832 2296 4288 5680
<< labels >>
flabel metal1 930 2354 1130 2538 0 FreeSans 800 0 0 0 vdd
port 2 nsew
flabel metal1 3676 246 3884 440 0 FreeSans 800 0 0 0 vss
port 4 nsew
flabel metal1 4582 2706 4856 2956 0 FreeSans 800 0 0 0 cp_bias
port 5 nsew
flabel metal1 20 1902 266 2174 0 FreeSans 800 0 0 0 ref
port 9 nsew
flabel metal3 5654 3087 5976 3409 0 FreeSans 800 0 0 0 out
port 7 nsew
<< end >>
