magic
tech sky130A
magscale 1 2
timestamp 1713428059
<< pwell >>
rect -386 -280 386 280
<< nmos >>
rect -200 -80 200 80
<< ndiff >>
rect -258 51 -200 80
rect -258 17 -246 51
rect -212 17 -200 51
rect -258 -17 -200 17
rect -258 -51 -246 -17
rect -212 -51 -200 -17
rect -258 -80 -200 -51
rect 200 51 258 80
rect 200 17 212 51
rect 246 17 258 51
rect 200 -17 258 17
rect 200 -51 212 -17
rect 246 -51 258 -17
rect 200 -80 258 -51
<< ndiffc >>
rect -246 17 -212 51
rect -246 -51 -212 -17
rect 212 17 246 51
rect 212 -51 246 -17
<< psubdiff >>
rect -360 220 -255 254
rect -221 220 -187 254
rect -153 220 -119 254
rect -85 220 -51 254
rect -17 220 17 254
rect 51 220 85 254
rect 119 220 153 254
rect 187 220 221 254
rect 255 220 360 254
rect -360 153 -326 220
rect -360 85 -326 119
rect 326 153 360 220
rect 326 85 360 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect 326 17 360 51
rect 326 -51 360 -17
rect -360 -119 -326 -85
rect -360 -220 -326 -153
rect 326 -119 360 -85
rect 326 -220 360 -153
rect -360 -254 -255 -220
rect -221 -254 -187 -220
rect -153 -254 -119 -220
rect -85 -254 -51 -220
rect -17 -254 17 -220
rect 51 -254 85 -220
rect 119 -254 153 -220
rect 187 -254 221 -220
rect 255 -254 360 -220
<< psubdiffcont >>
rect -255 220 -221 254
rect -187 220 -153 254
rect -119 220 -85 254
rect -51 220 -17 254
rect 17 220 51 254
rect 85 220 119 254
rect 153 220 187 254
rect 221 220 255 254
rect -360 119 -326 153
rect -360 51 -326 85
rect 326 119 360 153
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect 326 51 360 85
rect 326 -17 360 17
rect -360 -153 -326 -119
rect 326 -85 360 -51
rect 326 -153 360 -119
rect -255 -254 -221 -220
rect -187 -254 -153 -220
rect -119 -254 -85 -220
rect -51 -254 -17 -220
rect 17 -254 51 -220
rect 85 -254 119 -220
rect 153 -254 187 -220
rect 221 -254 255 -220
<< poly >>
rect -200 152 200 168
rect -200 118 -153 152
rect -119 118 -85 152
rect -51 118 -17 152
rect 17 118 51 152
rect 85 118 119 152
rect 153 118 200 152
rect -200 80 200 118
rect -200 -118 200 -80
rect -200 -152 -153 -118
rect -119 -152 -85 -118
rect -51 -152 -17 -118
rect 17 -152 51 -118
rect 85 -152 119 -118
rect 153 -152 200 -118
rect -200 -168 200 -152
<< polycont >>
rect -153 118 -119 152
rect -85 118 -51 152
rect -17 118 17 152
rect 51 118 85 152
rect 119 118 153 152
rect -153 -152 -119 -118
rect -85 -152 -51 -118
rect -17 -152 17 -118
rect 51 -152 85 -118
rect 119 -152 153 -118
<< locali >>
rect -360 220 -255 254
rect -221 220 -187 254
rect -153 220 -119 254
rect -85 220 -51 254
rect -17 220 17 254
rect 51 220 85 254
rect 119 220 153 254
rect 187 220 221 254
rect 255 220 360 254
rect -360 153 -326 220
rect 326 153 360 220
rect -360 85 -326 119
rect -200 118 -161 152
rect -119 118 -89 152
rect -51 118 -17 152
rect 17 118 51 152
rect 89 118 119 152
rect 161 118 200 152
rect 326 85 360 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -246 53 -212 84
rect -246 -17 -212 17
rect -246 -84 -212 -53
rect 212 53 246 84
rect 212 -17 246 17
rect 212 -84 246 -53
rect 326 17 360 51
rect 326 -51 360 -17
rect -360 -119 -326 -85
rect -200 -152 -161 -118
rect -119 -152 -89 -118
rect -51 -152 -17 -118
rect 17 -152 51 -118
rect 89 -152 119 -118
rect 161 -152 200 -118
rect 326 -119 360 -85
rect -360 -220 -326 -153
rect 326 -220 360 -153
rect -360 -254 -255 -220
rect -221 -254 -187 -220
rect -153 -254 -119 -220
rect -85 -254 -51 -220
rect -17 -254 17 -220
rect 51 -254 85 -220
rect 119 -254 153 -220
rect 187 -254 221 -220
rect 255 -254 360 -220
<< viali >>
rect -161 118 -153 152
rect -153 118 -127 152
rect -89 118 -85 152
rect -85 118 -55 152
rect -17 118 17 152
rect 55 118 85 152
rect 85 118 89 152
rect 127 118 153 152
rect 153 118 161 152
rect -246 51 -212 53
rect -246 19 -212 51
rect -246 -51 -212 -19
rect -246 -53 -212 -51
rect 212 51 246 53
rect 212 19 246 51
rect 212 -51 246 -19
rect 212 -53 246 -51
rect -161 -152 -153 -118
rect -153 -152 -127 -118
rect -89 -152 -85 -118
rect -85 -152 -55 -118
rect -17 -152 17 -118
rect 55 -152 85 -118
rect 85 -152 89 -118
rect 127 -152 153 -118
rect 153 -152 161 -118
<< metal1 >>
rect -196 152 196 158
rect -196 118 -161 152
rect -127 118 -89 152
rect -55 118 -17 152
rect 17 118 55 152
rect 89 118 127 152
rect 161 118 196 152
rect -196 112 196 118
rect -252 53 -206 80
rect -252 19 -246 53
rect -212 19 -206 53
rect -252 -19 -206 19
rect -252 -53 -246 -19
rect -212 -53 -206 -19
rect -252 -80 -206 -53
rect 206 53 252 80
rect 206 19 212 53
rect 246 19 252 53
rect 206 -19 252 19
rect 206 -53 212 -19
rect 246 -53 252 -19
rect 206 -80 252 -53
rect -196 -118 196 -112
rect -196 -152 -161 -118
rect -127 -152 -89 -118
rect -55 -152 -17 -118
rect 17 -152 55 -118
rect 89 -152 127 -118
rect 161 -152 196 -118
rect -196 -158 196 -152
<< properties >>
string FIXED_BBOX -342 -236 342 236
<< end >>
