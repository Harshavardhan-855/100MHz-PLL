magic
tech sky130A
magscale 1 2
timestamp 1709710021
<< error_s >>
rect 2692 1202 2974 1204
rect 2884 242 3018 244
rect 2912 214 2990 216
<< viali >>
rect 2524 -976 3220 -920
<< metal1 >>
rect 2688 1358 2938 2094
rect 2688 696 2698 1116
rect 2970 696 2980 1116
rect 3512 404 3522 630
rect 3736 404 3746 630
rect 2130 302 3326 304
rect 2112 242 3326 302
rect 2112 -158 2198 242
rect 2340 -98 2350 204
rect 2408 -98 2418 204
rect 2528 -92 2538 210
rect 2596 -92 2606 210
rect 2724 -92 2734 210
rect 2792 -92 2802 210
rect 2912 -86 2922 216
rect 2980 -86 2990 216
rect 3108 -94 3118 208
rect 3176 -94 3186 208
rect 3300 -96 3310 206
rect 3368 -96 3378 206
rect 1918 -358 2198 -158
rect 2112 -816 2198 -358
rect 2436 -768 2446 -482
rect 2508 -768 2518 -482
rect 2626 -766 2636 -480
rect 2698 -766 2708 -480
rect 2816 -770 2826 -484
rect 2888 -770 2898 -484
rect 3012 -772 3022 -486
rect 3084 -772 3094 -486
rect 3202 -774 3212 -488
rect 3274 -774 3284 -488
rect 2112 -868 3230 -816
rect 2132 -870 3230 -868
rect 2504 -998 2514 -904
rect 3278 -998 3288 -904
rect 2710 -1300 2720 -1058
rect 3026 -1300 3036 -1058
<< via1 >>
rect 2698 696 2970 1116
rect 3522 404 3736 630
rect 2350 -98 2408 204
rect 2538 -92 2596 210
rect 2734 -92 2792 210
rect 2922 -86 2980 216
rect 3118 -94 3176 208
rect 3310 -96 3368 206
rect 2446 -768 2508 -482
rect 2636 -766 2698 -480
rect 2826 -770 2888 -484
rect 3022 -772 3084 -486
rect 3212 -774 3274 -488
rect 2514 -920 3278 -904
rect 2514 -976 2524 -920
rect 2524 -976 3220 -920
rect 3220 -976 3278 -920
rect 2514 -998 3278 -976
rect 2720 -1300 3026 -1058
<< metal2 >>
rect 2698 1116 2970 1126
rect 2698 686 2970 696
rect 2700 650 2968 686
rect 2700 630 3744 650
rect 2700 404 3522 630
rect 3736 404 3744 630
rect 2700 392 3744 404
rect 2700 226 2968 392
rect 2350 204 2408 214
rect 2342 -84 2350 194
rect 2538 210 2596 220
rect 2408 -84 2538 194
rect 2350 -108 2408 -98
rect 2700 216 2980 226
rect 2700 210 2922 216
rect 2700 194 2734 210
rect 2596 -84 2734 194
rect 2538 -102 2596 -92
rect 2792 -84 2922 210
rect 2734 -102 2792 -92
rect 3118 208 3176 218
rect 2980 -84 3118 194
rect 2922 -96 2980 -86
rect 3310 206 3368 216
rect 3176 -84 3310 194
rect 3118 -104 3176 -94
rect 3368 -84 3370 194
rect 3310 -106 3368 -96
rect 2446 -482 2508 -472
rect 2440 -758 2446 -534
rect 2636 -480 2698 -470
rect 2508 -758 2636 -534
rect 2446 -778 2508 -768
rect 2826 -484 2888 -474
rect 2698 -758 2826 -534
rect 2636 -776 2698 -766
rect 2742 -770 2826 -758
rect 3022 -486 3084 -476
rect 2888 -758 3022 -534
rect 2888 -770 2978 -758
rect 2742 -894 2978 -770
rect 3212 -488 3274 -478
rect 3084 -758 3212 -534
rect 3022 -782 3084 -772
rect 3212 -784 3274 -774
rect 2514 -904 3278 -894
rect 2514 -1008 3278 -998
rect 2742 -1048 2978 -1008
rect 2720 -1058 3026 -1048
rect 2720 -1310 3026 -1300
use sky130_fd_pr__nfet_01v8_P4JNYZ  XM1
timestamp 1709710021
transform 1 0 2859 0 1 -288
box -647 -710 647 710
use sky130_fd_pr__res_high_po_1p41_DQDBL4  XR1
timestamp 1709710021
transform -1 0 2833 0 1 1168
box -307 -632 307 632
<< labels >>
flabel metal1 1918 -358 2118 -158 0 FreeSans 256 0 0 0 inp
port 2 nsew
flabel via1 2768 -1292 2968 -1092 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 2692 1874 2892 2074 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel via1 3532 412 3732 612 0 FreeSans 256 0 0 0 out
port 1 nsew
<< end >>
