magic
tech sky130A
magscale 1 2
timestamp 1709710021
<< error_p >>
rect -365 5072 -307 5078
rect -173 5072 -115 5078
rect 19 5072 77 5078
rect 211 5072 269 5078
rect 403 5072 461 5078
rect -365 5038 -353 5072
rect -173 5038 -161 5072
rect 19 5038 31 5072
rect 211 5038 223 5072
rect 403 5038 415 5072
rect -365 5032 -307 5038
rect -173 5032 -115 5038
rect 19 5032 77 5038
rect 211 5032 269 5038
rect 403 5032 461 5038
rect -461 -5038 -403 -5032
rect -269 -5038 -211 -5032
rect -77 -5038 -19 -5032
rect 115 -5038 173 -5032
rect 307 -5038 365 -5032
rect -461 -5072 -449 -5038
rect -269 -5072 -257 -5038
rect -77 -5072 -65 -5038
rect 115 -5072 127 -5038
rect 307 -5072 319 -5038
rect -461 -5078 -403 -5072
rect -269 -5078 -211 -5072
rect -77 -5078 -19 -5072
rect 115 -5078 173 -5072
rect 307 -5078 365 -5072
<< pwell >>
rect -647 -5210 647 5210
<< nmos >>
rect -447 -5000 -417 5000
rect -351 -5000 -321 5000
rect -255 -5000 -225 5000
rect -159 -5000 -129 5000
rect -63 -5000 -33 5000
rect 33 -5000 63 5000
rect 129 -5000 159 5000
rect 225 -5000 255 5000
rect 321 -5000 351 5000
rect 417 -5000 447 5000
<< ndiff >>
rect -509 4988 -447 5000
rect -509 -4988 -497 4988
rect -463 -4988 -447 4988
rect -509 -5000 -447 -4988
rect -417 4988 -351 5000
rect -417 -4988 -401 4988
rect -367 -4988 -351 4988
rect -417 -5000 -351 -4988
rect -321 4988 -255 5000
rect -321 -4988 -305 4988
rect -271 -4988 -255 4988
rect -321 -5000 -255 -4988
rect -225 4988 -159 5000
rect -225 -4988 -209 4988
rect -175 -4988 -159 4988
rect -225 -5000 -159 -4988
rect -129 4988 -63 5000
rect -129 -4988 -113 4988
rect -79 -4988 -63 4988
rect -129 -5000 -63 -4988
rect -33 4988 33 5000
rect -33 -4988 -17 4988
rect 17 -4988 33 4988
rect -33 -5000 33 -4988
rect 63 4988 129 5000
rect 63 -4988 79 4988
rect 113 -4988 129 4988
rect 63 -5000 129 -4988
rect 159 4988 225 5000
rect 159 -4988 175 4988
rect 209 -4988 225 4988
rect 159 -5000 225 -4988
rect 255 4988 321 5000
rect 255 -4988 271 4988
rect 305 -4988 321 4988
rect 255 -5000 321 -4988
rect 351 4988 417 5000
rect 351 -4988 367 4988
rect 401 -4988 417 4988
rect 351 -5000 417 -4988
rect 447 4988 509 5000
rect 447 -4988 463 4988
rect 497 -4988 509 4988
rect 447 -5000 509 -4988
<< ndiffc >>
rect -497 -4988 -463 4988
rect -401 -4988 -367 4988
rect -305 -4988 -271 4988
rect -209 -4988 -175 4988
rect -113 -4988 -79 4988
rect -17 -4988 17 4988
rect 79 -4988 113 4988
rect 175 -4988 209 4988
rect 271 -4988 305 4988
rect 367 -4988 401 4988
rect 463 -4988 497 4988
<< psubdiff >>
rect -611 5140 -515 5174
rect 515 5140 611 5174
rect -611 5078 -577 5140
rect 577 5078 611 5140
rect -611 -5140 -577 -5078
rect 577 -5140 611 -5078
rect -611 -5174 -515 -5140
rect 515 -5174 611 -5140
<< psubdiffcont >>
rect -515 5140 515 5174
rect -611 -5078 -577 5078
rect 577 -5078 611 5078
rect -515 -5174 515 -5140
<< poly >>
rect -369 5072 -303 5088
rect -369 5038 -353 5072
rect -319 5038 -303 5072
rect -447 5000 -417 5026
rect -369 5022 -303 5038
rect -177 5072 -111 5088
rect -177 5038 -161 5072
rect -127 5038 -111 5072
rect -351 5000 -321 5022
rect -255 5000 -225 5026
rect -177 5022 -111 5038
rect 15 5072 81 5088
rect 15 5038 31 5072
rect 65 5038 81 5072
rect -159 5000 -129 5022
rect -63 5000 -33 5026
rect 15 5022 81 5038
rect 207 5072 273 5088
rect 207 5038 223 5072
rect 257 5038 273 5072
rect 33 5000 63 5022
rect 129 5000 159 5026
rect 207 5022 273 5038
rect 399 5072 465 5088
rect 399 5038 415 5072
rect 449 5038 465 5072
rect 225 5000 255 5022
rect 321 5000 351 5026
rect 399 5022 465 5038
rect 417 5000 447 5022
rect -447 -5022 -417 -5000
rect -465 -5038 -399 -5022
rect -351 -5026 -321 -5000
rect -255 -5022 -225 -5000
rect -465 -5072 -449 -5038
rect -415 -5072 -399 -5038
rect -465 -5088 -399 -5072
rect -273 -5038 -207 -5022
rect -159 -5026 -129 -5000
rect -63 -5022 -33 -5000
rect -273 -5072 -257 -5038
rect -223 -5072 -207 -5038
rect -273 -5088 -207 -5072
rect -81 -5038 -15 -5022
rect 33 -5026 63 -5000
rect 129 -5022 159 -5000
rect -81 -5072 -65 -5038
rect -31 -5072 -15 -5038
rect -81 -5088 -15 -5072
rect 111 -5038 177 -5022
rect 225 -5026 255 -5000
rect 321 -5022 351 -5000
rect 111 -5072 127 -5038
rect 161 -5072 177 -5038
rect 111 -5088 177 -5072
rect 303 -5038 369 -5022
rect 417 -5026 447 -5000
rect 303 -5072 319 -5038
rect 353 -5072 369 -5038
rect 303 -5088 369 -5072
<< polycont >>
rect -353 5038 -319 5072
rect -161 5038 -127 5072
rect 31 5038 65 5072
rect 223 5038 257 5072
rect 415 5038 449 5072
rect -449 -5072 -415 -5038
rect -257 -5072 -223 -5038
rect -65 -5072 -31 -5038
rect 127 -5072 161 -5038
rect 319 -5072 353 -5038
<< locali >>
rect -611 5140 -515 5174
rect 515 5140 611 5174
rect -611 5078 -577 5140
rect 577 5078 611 5140
rect -369 5038 -353 5072
rect -319 5038 -303 5072
rect -177 5038 -161 5072
rect -127 5038 -111 5072
rect 15 5038 31 5072
rect 65 5038 81 5072
rect 207 5038 223 5072
rect 257 5038 273 5072
rect 399 5038 415 5072
rect 449 5038 465 5072
rect -497 4988 -463 5004
rect -497 -5004 -463 -4988
rect -401 4988 -367 5004
rect -401 -5004 -367 -4988
rect -305 4988 -271 5004
rect -305 -5004 -271 -4988
rect -209 4988 -175 5004
rect -209 -5004 -175 -4988
rect -113 4988 -79 5004
rect -113 -5004 -79 -4988
rect -17 4988 17 5004
rect -17 -5004 17 -4988
rect 79 4988 113 5004
rect 79 -5004 113 -4988
rect 175 4988 209 5004
rect 175 -5004 209 -4988
rect 271 4988 305 5004
rect 271 -5004 305 -4988
rect 367 4988 401 5004
rect 367 -5004 401 -4988
rect 463 4988 497 5004
rect 463 -5004 497 -4988
rect -465 -5072 -449 -5038
rect -415 -5072 -399 -5038
rect -273 -5072 -257 -5038
rect -223 -5072 -207 -5038
rect -81 -5072 -65 -5038
rect -31 -5072 -15 -5038
rect 111 -5072 127 -5038
rect 161 -5072 177 -5038
rect 303 -5072 319 -5038
rect 353 -5072 369 -5038
rect -611 -5140 -577 -5078
rect 577 -5140 611 -5078
rect -611 -5174 -515 -5140
rect 515 -5174 611 -5140
<< viali >>
rect -353 5038 -319 5072
rect -161 5038 -127 5072
rect 31 5038 65 5072
rect 223 5038 257 5072
rect 415 5038 449 5072
rect -497 -4988 -463 4988
rect -401 -4988 -367 4988
rect -305 -4988 -271 4988
rect -209 -4988 -175 4988
rect -113 -4988 -79 4988
rect -17 -4988 17 4988
rect 79 -4988 113 4988
rect 175 -4988 209 4988
rect 271 -4988 305 4988
rect 367 -4988 401 4988
rect 463 -4988 497 4988
rect -449 -5072 -415 -5038
rect -257 -5072 -223 -5038
rect -65 -5072 -31 -5038
rect 127 -5072 161 -5038
rect 319 -5072 353 -5038
<< metal1 >>
rect -365 5072 -307 5078
rect -365 5038 -353 5072
rect -319 5038 -307 5072
rect -365 5032 -307 5038
rect -173 5072 -115 5078
rect -173 5038 -161 5072
rect -127 5038 -115 5072
rect -173 5032 -115 5038
rect 19 5072 77 5078
rect 19 5038 31 5072
rect 65 5038 77 5072
rect 19 5032 77 5038
rect 211 5072 269 5078
rect 211 5038 223 5072
rect 257 5038 269 5072
rect 211 5032 269 5038
rect 403 5072 461 5078
rect 403 5038 415 5072
rect 449 5038 461 5072
rect 403 5032 461 5038
rect -503 4988 -457 5000
rect -503 -4988 -497 4988
rect -463 -4988 -457 4988
rect -503 -5000 -457 -4988
rect -407 4988 -361 5000
rect -407 -4988 -401 4988
rect -367 -4988 -361 4988
rect -407 -5000 -361 -4988
rect -311 4988 -265 5000
rect -311 -4988 -305 4988
rect -271 -4988 -265 4988
rect -311 -5000 -265 -4988
rect -215 4988 -169 5000
rect -215 -4988 -209 4988
rect -175 -4988 -169 4988
rect -215 -5000 -169 -4988
rect -119 4988 -73 5000
rect -119 -4988 -113 4988
rect -79 -4988 -73 4988
rect -119 -5000 -73 -4988
rect -23 4988 23 5000
rect -23 -4988 -17 4988
rect 17 -4988 23 4988
rect -23 -5000 23 -4988
rect 73 4988 119 5000
rect 73 -4988 79 4988
rect 113 -4988 119 4988
rect 73 -5000 119 -4988
rect 169 4988 215 5000
rect 169 -4988 175 4988
rect 209 -4988 215 4988
rect 169 -5000 215 -4988
rect 265 4988 311 5000
rect 265 -4988 271 4988
rect 305 -4988 311 4988
rect 265 -5000 311 -4988
rect 361 4988 407 5000
rect 361 -4988 367 4988
rect 401 -4988 407 4988
rect 361 -5000 407 -4988
rect 457 4988 503 5000
rect 457 -4988 463 4988
rect 497 -4988 503 4988
rect 457 -5000 503 -4988
rect -461 -5038 -403 -5032
rect -461 -5072 -449 -5038
rect -415 -5072 -403 -5038
rect -461 -5078 -403 -5072
rect -269 -5038 -211 -5032
rect -269 -5072 -257 -5038
rect -223 -5072 -211 -5038
rect -269 -5078 -211 -5072
rect -77 -5038 -19 -5032
rect -77 -5072 -65 -5038
rect -31 -5072 -19 -5038
rect -77 -5078 -19 -5072
rect 115 -5038 173 -5032
rect 115 -5072 127 -5038
rect 161 -5072 173 -5038
rect 115 -5078 173 -5072
rect 307 -5038 365 -5032
rect 307 -5072 319 -5038
rect 353 -5072 365 -5038
rect 307 -5078 365 -5072
<< properties >>
string FIXED_BBOX -594 -5157 594 5157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 50.0 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
