magic
tech sky130A
magscale 1 2
timestamp 1709710021
<< error_p >>
rect -365 572 -307 578
rect -173 572 -115 578
rect 19 572 77 578
rect 211 572 269 578
rect 403 572 461 578
rect -365 538 -353 572
rect -173 538 -161 572
rect 19 538 31 572
rect 211 538 223 572
rect 403 538 415 572
rect -365 532 -307 538
rect -173 532 -115 538
rect 19 532 77 538
rect 211 532 269 538
rect 403 532 461 538
rect -461 -538 -403 -532
rect -269 -538 -211 -532
rect -77 -538 -19 -532
rect 115 -538 173 -532
rect 307 -538 365 -532
rect -461 -572 -449 -538
rect -269 -572 -257 -538
rect -77 -572 -65 -538
rect 115 -572 127 -538
rect 307 -572 319 -538
rect -461 -578 -403 -572
rect -269 -578 -211 -572
rect -77 -578 -19 -572
rect 115 -578 173 -572
rect 307 -578 365 -572
<< pwell >>
rect -647 -710 647 710
<< nmos >>
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
<< ndiff >>
rect -509 488 -447 500
rect -509 -488 -497 488
rect -463 -488 -447 488
rect -509 -500 -447 -488
rect -417 488 -351 500
rect -417 -488 -401 488
rect -367 -488 -351 488
rect -417 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 417 500
rect 351 -488 367 488
rect 401 -488 417 488
rect 351 -500 417 -488
rect 447 488 509 500
rect 447 -488 463 488
rect 497 -488 509 488
rect 447 -500 509 -488
<< ndiffc >>
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
<< psubdiff >>
rect -611 640 -515 674
rect 515 640 611 674
rect -611 578 -577 640
rect 577 578 611 640
rect -611 -640 -577 -578
rect 577 -640 611 -578
rect -611 -674 -515 -640
rect 515 -674 611 -640
<< psubdiffcont >>
rect -515 640 515 674
rect -611 -578 -577 578
rect 577 -578 611 578
rect -515 -674 515 -640
<< poly >>
rect -369 572 -303 588
rect -369 538 -353 572
rect -319 538 -303 572
rect -447 500 -417 526
rect -369 522 -303 538
rect -177 572 -111 588
rect -177 538 -161 572
rect -127 538 -111 572
rect -351 500 -321 522
rect -255 500 -225 526
rect -177 522 -111 538
rect 15 572 81 588
rect 15 538 31 572
rect 65 538 81 572
rect -159 500 -129 522
rect -63 500 -33 526
rect 15 522 81 538
rect 207 572 273 588
rect 207 538 223 572
rect 257 538 273 572
rect 33 500 63 522
rect 129 500 159 526
rect 207 522 273 538
rect 399 572 465 588
rect 399 538 415 572
rect 449 538 465 572
rect 225 500 255 522
rect 321 500 351 526
rect 399 522 465 538
rect 417 500 447 522
rect -447 -522 -417 -500
rect -465 -538 -399 -522
rect -351 -526 -321 -500
rect -255 -522 -225 -500
rect -465 -572 -449 -538
rect -415 -572 -399 -538
rect -465 -588 -399 -572
rect -273 -538 -207 -522
rect -159 -526 -129 -500
rect -63 -522 -33 -500
rect -273 -572 -257 -538
rect -223 -572 -207 -538
rect -273 -588 -207 -572
rect -81 -538 -15 -522
rect 33 -526 63 -500
rect 129 -522 159 -500
rect -81 -572 -65 -538
rect -31 -572 -15 -538
rect -81 -588 -15 -572
rect 111 -538 177 -522
rect 225 -526 255 -500
rect 321 -522 351 -500
rect 111 -572 127 -538
rect 161 -572 177 -538
rect 111 -588 177 -572
rect 303 -538 369 -522
rect 417 -526 447 -500
rect 303 -572 319 -538
rect 353 -572 369 -538
rect 303 -588 369 -572
<< polycont >>
rect -353 538 -319 572
rect -161 538 -127 572
rect 31 538 65 572
rect 223 538 257 572
rect 415 538 449 572
rect -449 -572 -415 -538
rect -257 -572 -223 -538
rect -65 -572 -31 -538
rect 127 -572 161 -538
rect 319 -572 353 -538
<< locali >>
rect -611 640 -515 674
rect 515 640 611 674
rect -611 578 -577 640
rect 577 578 611 640
rect -369 538 -353 572
rect -319 538 -303 572
rect -177 538 -161 572
rect -127 538 -111 572
rect 15 538 31 572
rect 65 538 81 572
rect 207 538 223 572
rect 257 538 273 572
rect 399 538 415 572
rect 449 538 465 572
rect -497 488 -463 504
rect -497 -504 -463 -488
rect -401 488 -367 504
rect -401 -504 -367 -488
rect -305 488 -271 504
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect 271 488 305 504
rect 271 -504 305 -488
rect 367 488 401 504
rect 367 -504 401 -488
rect 463 488 497 504
rect 463 -504 497 -488
rect -465 -572 -449 -538
rect -415 -572 -399 -538
rect -273 -572 -257 -538
rect -223 -572 -207 -538
rect -81 -572 -65 -538
rect -31 -572 -15 -538
rect 111 -572 127 -538
rect 161 -572 177 -538
rect 303 -572 319 -538
rect 353 -572 369 -538
rect -611 -640 -577 -578
rect 577 -640 611 -578
rect -611 -674 -515 -640
rect 515 -674 611 -640
<< viali >>
rect -353 538 -319 572
rect -161 538 -127 572
rect 31 538 65 572
rect 223 538 257 572
rect 415 538 449 572
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect -449 -572 -415 -538
rect -257 -572 -223 -538
rect -65 -572 -31 -538
rect 127 -572 161 -538
rect 319 -572 353 -538
<< metal1 >>
rect -365 572 -307 578
rect -365 538 -353 572
rect -319 538 -307 572
rect -365 532 -307 538
rect -173 572 -115 578
rect -173 538 -161 572
rect -127 538 -115 572
rect -173 532 -115 538
rect 19 572 77 578
rect 19 538 31 572
rect 65 538 77 572
rect 19 532 77 538
rect 211 572 269 578
rect 211 538 223 572
rect 257 538 269 572
rect 211 532 269 538
rect 403 572 461 578
rect 403 538 415 572
rect 449 538 461 572
rect 403 532 461 538
rect -503 488 -457 500
rect -503 -488 -497 488
rect -463 -488 -457 488
rect -503 -500 -457 -488
rect -407 488 -361 500
rect -407 -488 -401 488
rect -367 -488 -361 488
rect -407 -500 -361 -488
rect -311 488 -265 500
rect -311 -488 -305 488
rect -271 -488 -265 488
rect -311 -500 -265 -488
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect 265 488 311 500
rect 265 -488 271 488
rect 305 -488 311 488
rect 265 -500 311 -488
rect 361 488 407 500
rect 361 -488 367 488
rect 401 -488 407 488
rect 361 -500 407 -488
rect 457 488 503 500
rect 457 -488 463 488
rect 497 -488 503 488
rect 457 -500 503 -488
rect -461 -538 -403 -532
rect -461 -572 -449 -538
rect -415 -572 -403 -538
rect -461 -578 -403 -572
rect -269 -538 -211 -532
rect -269 -572 -257 -538
rect -223 -572 -211 -538
rect -269 -578 -211 -572
rect -77 -538 -19 -532
rect -77 -572 -65 -538
rect -31 -572 -19 -538
rect -77 -578 -19 -572
rect 115 -538 173 -532
rect 115 -572 127 -538
rect 161 -572 173 -538
rect 115 -578 173 -572
rect 307 -538 365 -532
rect 307 -572 319 -538
rect 353 -572 365 -538
rect 307 -578 365 -572
<< properties >>
string FIXED_BBOX -594 -657 594 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
