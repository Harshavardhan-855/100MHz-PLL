* NGSPICE file created from cs.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_1p41_DQDBL4 a_n141_n466# a_n271_n596# a_n141_34#
X0 a_n141_34# a_n141_n466# a_n271_n596# sky130_fd_pr__res_high_po_1p41 l=0.5
C0 a_n141_n466# a_n141_34# 0.168219f
C1 a_n141_n466# a_n271_n596# 0.744526f
C2 a_n141_34# a_n271_n596# 0.744526f
.ends

.subckt sky130_fd_pr__nfet_01v8_P4JNYZ a_n129_n500# a_n81_n588# a_63_n500# a_n177_522#
+ a_n225_n500# a_n321_n500# a_n369_522# a_n33_n500# a_n509_n500# a_303_n588# a_447_n500#
+ a_n465_n588# a_399_522# a_159_n500# a_111_n588# a_15_522# a_n273_n588# a_255_n500#
+ a_n611_n674# a_207_522# a_351_n500# a_n417_n500#
X0 a_n417_n500# a_n465_n588# a_n509_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X1 a_n33_n500# a_n81_n588# a_n129_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X2 a_351_n500# a_303_n588# a_255_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X3 a_255_n500# a_207_522# a_159_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X4 a_n321_n500# a_n369_522# a_n417_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X5 a_159_n500# a_111_n588# a_63_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X6 a_n225_n500# a_n273_n588# a_n321_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X7 a_447_n500# a_399_522# a_351_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X8 a_63_n500# a_15_522# a_n33_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X9 a_n129_n500# a_n177_522# a_n225_n500# a_n611_n674# sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
C0 a_n273_n588# a_n225_n500# 0.029899f
C1 a_n177_522# a_n369_522# 0.02473f
C2 a_n33_n500# a_n129_n500# 0.735411f
C3 a_207_522# a_159_n500# 0.029899f
C4 a_n33_n500# a_63_n500# 0.735411f
C5 a_n273_n588# a_n81_n588# 0.02473f
C6 a_399_522# a_207_522# 0.02473f
C7 a_n273_n588# a_n177_522# 0.013333f
C8 a_15_522# a_n81_n588# 0.013333f
C9 a_n321_n500# a_n369_522# 0.029899f
C10 a_15_522# a_n177_522# 0.02473f
C11 a_303_n588# a_111_n588# 0.02473f
C12 a_111_n588# a_n81_n588# 0.02473f
C13 a_351_n500# a_255_n500# 0.735411f
C14 a_n509_n500# a_n465_n588# 0.029899f
C15 a_n321_n500# a_n273_n588# 0.029899f
C16 a_399_522# a_447_n500# 0.029899f
C17 a_15_522# a_n33_n500# 0.029899f
C18 a_n369_522# a_n465_n588# 0.013333f
C19 a_399_522# a_303_n588# 0.013333f
C20 a_n321_n500# a_n417_n500# 0.735411f
C21 a_207_522# a_303_n588# 0.013333f
C22 a_n273_n588# a_n465_n588# 0.02473f
C23 a_n273_n588# a_n369_522# 0.013333f
C24 a_15_522# a_63_n500# 0.029899f
C25 a_n509_n500# a_n417_n500# 0.735411f
C26 a_n417_n500# a_n465_n588# 0.029899f
C27 a_63_n500# a_111_n588# 0.029899f
C28 a_n225_n500# a_n177_522# 0.029899f
C29 a_n417_n500# a_n369_522# 0.029899f
C30 a_399_522# a_351_n500# 0.029899f
C31 a_n81_n588# a_n177_522# 0.013333f
C32 a_63_n500# a_159_n500# 0.735411f
C33 a_159_n500# a_255_n500# 0.735411f
C34 a_n321_n500# a_n225_n500# 0.735411f
C35 a_15_522# a_111_n588# 0.013333f
C36 a_207_522# a_255_n500# 0.029899f
C37 a_n33_n500# a_n81_n588# 0.029899f
C38 a_351_n500# a_447_n500# 0.735411f
C39 a_n225_n500# a_n129_n500# 0.735411f
C40 a_351_n500# a_303_n588# 0.029899f
C41 a_159_n500# a_111_n588# 0.029899f
C42 a_15_522# a_207_522# 0.02473f
C43 a_n129_n500# a_n81_n588# 0.029899f
C44 a_n129_n500# a_n177_522# 0.029899f
C45 a_303_n588# a_255_n500# 0.029899f
C46 a_207_522# a_111_n588# 0.013333f
C47 a_447_n500# a_n611_n674# 0.544674f
C48 a_351_n500# a_n611_n674# 0.073056f
C49 a_255_n500# a_n611_n674# 0.073056f
C50 a_159_n500# a_n611_n674# 0.073056f
C51 a_63_n500# a_n611_n674# 0.073056f
C52 a_n33_n500# a_n611_n674# 0.073056f
C53 a_n129_n500# a_n611_n674# 0.073056f
C54 a_n225_n500# a_n611_n674# 0.073056f
C55 a_n321_n500# a_n611_n674# 0.073056f
C56 a_n417_n500# a_n611_n674# 0.073056f
C57 a_n509_n500# a_n611_n674# 0.544674f
C58 a_303_n588# a_n611_n674# 0.170156f
C59 a_399_522# a_n611_n674# 0.182024f
C60 a_111_n588# a_n611_n674# 0.150661f
C61 a_207_522# a_n611_n674# 0.150691f
C62 a_n81_n588# a_n611_n674# 0.150649f
C63 a_15_522# a_n611_n674# 0.150649f
C64 a_n273_n588# a_n611_n674# 0.150691f
C65 a_n177_522# a_n611_n674# 0.150661f
C66 a_n465_n588# a_n611_n674# 0.182024f
C67 a_n369_522# a_n611_n674# 0.170156f
.ends

.subckt cs_pex vdd out inp vss
XXR1 out vss vdd sky130_fd_pr__res_high_po_1p41_DQDBL4
XXM1 out inp out inp vss out inp vss out inp out inp inp vss inp inp inp out vss inp
+ vss vss sky130_fd_pr__nfet_01v8_P4JNYZ
C0 vdd inp 6.41e-19
C1 vdd out 0.042142f
C2 inp out 1.056944f
C3 inp vss 3.454313f
C4 out vss 4.496978f
C5 vdd vss 1.04611f
.ends

