magic
tech sky130A
timestamp 1711524713
<< metal4 >>
rect 200 22476 230 22576
rect 568 22476 598 22576
rect 936 22476 966 22576
rect 1304 22476 1334 22576
rect 1672 22476 1702 22576
rect 2040 22476 2070 22576
rect 2408 22476 2438 22576
rect 2776 22476 2806 22576
rect 3144 22476 3174 22576
rect 3512 22476 3542 22576
rect 3880 22476 3910 22576
rect 4248 22476 4278 22576
rect 4616 22476 4646 22576
rect 4984 22476 5014 22576
rect 5352 22476 5382 22576
rect 5720 22476 5750 22576
rect 6088 22476 6118 22576
rect 6456 22476 6486 22576
rect 6824 22476 6854 22576
rect 7192 22476 7222 22576
rect 7560 22476 7590 22576
rect 7928 22476 7958 22576
rect 8296 22476 8326 22576
rect 8664 22476 8694 22576
rect 9032 22476 9062 22576
rect 9400 22476 9430 22576
rect 9768 22476 9798 22576
rect 10136 22476 10166 22576
rect 10504 22476 10534 22576
rect 10872 22476 10902 22576
rect 11240 22476 11270 22576
rect 11608 22476 11638 22576
rect 11976 22476 12006 22576
rect 12344 22476 12374 22576
rect 12712 22476 12742 22576
rect 13080 22476 13110 22576
rect 13448 22476 13478 22576
rect 13816 22476 13846 22576
rect 14184 22476 14214 22576
rect 14552 22476 14582 22576
rect 14920 22476 14950 22576
rect 15288 22476 15318 22576
rect 15656 22476 15686 22576
rect 369 0 429 100
rect 2577 0 2637 100
rect 4785 0 4845 100
rect 6993 0 7053 100
rect 9201 0 9261 100
rect 11409 0 11469 100
rect 13617 0 13677 100
rect 15825 0 15885 100
<< labels >>
flabel metal4 s 568 22476 598 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 200 22476 230 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 936 22476 966 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 369 0 429 100 0 FreeSans 480 180 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 2577 0 2637 100 0 FreeSans 480 180 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 4785 0 4845 100 0 FreeSans 480 180 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 6993 0 7053 100 0 FreeSans 480 180 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 9201 0 9261 100 0 FreeSans 480 180 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11409 0 11469 100 0 FreeSans 480 180 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 13617 0 13677 100 0 FreeSans 480 180 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 15825 0 15885 100 0 FreeSans 480 180 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 1304 22476 1334 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 1672 22476 1702 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 2040 22476 2070 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 2408 22476 2438 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 2776 22476 2806 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 3144 22476 3174 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 3512 22476 3542 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 3880 22476 3910 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 4248 22476 4278 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 4616 22476 4646 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 4984 22476 5014 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 5352 22476 5382 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 5720 22476 5750 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 6088 22476 6118 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 6456 22476 6486 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 6824 22476 6854 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 13080 22476 13110 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 13448 22476 13478 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 13816 22476 13846 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 14184 22476 14214 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 14552 22476 14582 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 14920 22476 14950 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 15288 22476 15318 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 15656 22476 15686 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 10136 22476 10166 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10504 22476 10534 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10872 22476 10902 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 11240 22476 11270 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 11608 22476 11638 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11976 22476 12006 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 12344 22476 12374 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 12712 22476 12742 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 7192 22476 7222 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 7560 22476 7590 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 7928 22476 7958 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8296 22476 8326 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8664 22476 8694 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 9032 22476 9062 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 9400 22476 9430 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 9768 22476 9798 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 50876 22576
<< end >>
