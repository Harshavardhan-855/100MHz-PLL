magic
tech sky130A
magscale 1 2
timestamp 1713418708
<< checkpaint >>
rect -1313 -114 1629 45
rect -1313 -220 2796 -114
rect -1313 -326 3564 -220
rect -1313 -3313 4332 -326
rect -146 -3472 4332 -3313
rect 622 -3578 4332 -3472
rect 1390 -3684 4332 -3578
<< error_s >>
rect 129 -1353 187 -1347
rect 129 -1372 141 -1353
rect 129 -1393 187 -1372
rect 101 -1421 200 -1400
rect 299 -1486 333 -1468
rect 299 -1522 369 -1486
rect 1296 -1512 1354 -1506
rect 316 -1556 387 -1522
rect 697 -1556 732 -1522
rect 1150 -1539 1184 -1521
rect 316 -2017 386 -1556
rect 698 -1575 732 -1556
rect 513 -1624 571 -1618
rect 513 -1658 525 -1624
rect 513 -1664 571 -1658
rect 513 -1934 571 -1928
rect 513 -1968 525 -1934
rect 513 -1974 571 -1968
rect 316 -2053 369 -2017
rect 717 -2070 732 -1575
rect 751 -1609 786 -1575
rect 751 -2070 785 -1609
rect 912 -1677 970 -1671
rect 912 -1711 924 -1677
rect 912 -1717 970 -1711
rect 912 -1987 970 -1981
rect 912 -2021 924 -1987
rect 912 -2027 970 -2021
rect 751 -2104 766 -2070
rect 1114 -2123 1184 -1539
rect 1296 -1546 1308 -1512
rect 1296 -1552 1354 -1546
rect 2064 -1618 2122 -1612
rect 1466 -1645 1500 -1627
rect 1918 -1645 1952 -1627
rect 1466 -1681 1536 -1645
rect 1483 -1715 1554 -1681
rect 1296 -2040 1354 -2034
rect 1296 -2074 1308 -2040
rect 1296 -2080 1354 -2074
rect 1114 -2159 1167 -2123
rect 1483 -2176 1553 -1715
rect 1680 -1783 1738 -1777
rect 1680 -1817 1692 -1783
rect 1680 -1823 1738 -1817
rect 1680 -2093 1738 -2087
rect 1680 -2127 1692 -2093
rect 1680 -2133 1738 -2127
rect 1483 -2212 1536 -2176
rect 1882 -2229 1952 -1645
rect 2064 -1652 2076 -1618
rect 2064 -1658 2122 -1652
rect 2234 -1751 2268 -1733
rect 2234 -1787 2304 -1751
rect 2251 -1821 2322 -1787
rect 2064 -2146 2122 -2140
rect 2064 -2180 2076 -2146
rect 2064 -2186 2122 -2180
rect 1882 -2265 1935 -2229
rect 2251 -2282 2321 -1821
rect 2448 -1889 2506 -1883
rect 2448 -1923 2460 -1889
rect 2448 -1929 2506 -1923
rect 2448 -2199 2506 -2193
rect 2448 -2233 2460 -2199
rect 2448 -2239 2506 -2233
rect 2251 -2318 2304 -2282
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__pfet_01v8_XGAKDL  XM1
timestamp 0
transform 1 0 158 0 1 -1634
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_PSFW3M  XM2
timestamp 0
transform 1 0 542 0 1 -1796
box -226 -310 226 310
use sky130_fd_pr__nfet_01v8_PSFW3M  XM3
timestamp 0
transform 1 0 941 0 1 -1849
box -226 -310 226 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XM4
timestamp 0
transform 1 0 1325 0 1 -1793
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_PSFW3M  XM5
timestamp 0
transform 1 0 1709 0 1 -1955
box -226 -310 226 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XM6
timestamp 0
transform 1 0 2093 0 1 -1899
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_PSFW3M  XM7
timestamp 0
transform 1 0 2477 0 1 -2061
box -226 -310 226 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XM8
timestamp 0
transform 1 0 2861 0 1 -2005
box -211 -419 211 419
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 qa
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 cp_out
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 qb
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 cp_bias
port 5 nsew
<< end >>
