magic
tech sky130A
magscale 1 2
timestamp 1713432778
<< metal3 >>
rect -9378 8972 -3286 9000
rect -9378 3188 -3370 8972
rect -3306 3188 -3286 8972
rect -9378 3160 -3286 3188
rect -3046 8972 3046 9000
rect -3046 3188 2962 8972
rect 3026 3188 3046 8972
rect -3046 3160 3046 3188
rect 3286 8972 9378 9000
rect 3286 3188 9294 8972
rect 9358 3188 9378 8972
rect 3286 3160 9378 3188
rect -9378 2892 -3286 2920
rect -9378 -2892 -3370 2892
rect -3306 -2892 -3286 2892
rect -9378 -2920 -3286 -2892
rect -3046 2892 3046 2920
rect -3046 -2892 2962 2892
rect 3026 -2892 3046 2892
rect -3046 -2920 3046 -2892
rect 3286 2892 9378 2920
rect 3286 -2892 9294 2892
rect 9358 -2892 9378 2892
rect 3286 -2920 9378 -2892
rect -9378 -3188 -3286 -3160
rect -9378 -8972 -3370 -3188
rect -3306 -8972 -3286 -3188
rect -9378 -9000 -3286 -8972
rect -3046 -3188 3046 -3160
rect -3046 -8972 2962 -3188
rect 3026 -8972 3046 -3188
rect -3046 -9000 3046 -8972
rect 3286 -3188 9378 -3160
rect 3286 -8972 9294 -3188
rect 9358 -8972 9378 -3188
rect 3286 -9000 9378 -8972
<< via3 >>
rect -3370 3188 -3306 8972
rect 2962 3188 3026 8972
rect 9294 3188 9358 8972
rect -3370 -2892 -3306 2892
rect 2962 -2892 3026 2892
rect 9294 -2892 9358 2892
rect -3370 -8972 -3306 -3188
rect 2962 -8972 3026 -3188
rect 9294 -8972 9358 -3188
<< mimcap >>
rect -9338 8920 -3618 8960
rect -9338 3240 -9298 8920
rect -3658 3240 -3618 8920
rect -9338 3200 -3618 3240
rect -3006 8920 2714 8960
rect -3006 3240 -2966 8920
rect 2674 3240 2714 8920
rect -3006 3200 2714 3240
rect 3326 8920 9046 8960
rect 3326 3240 3366 8920
rect 9006 3240 9046 8920
rect 3326 3200 9046 3240
rect -9338 2840 -3618 2880
rect -9338 -2840 -9298 2840
rect -3658 -2840 -3618 2840
rect -9338 -2880 -3618 -2840
rect -3006 2840 2714 2880
rect -3006 -2840 -2966 2840
rect 2674 -2840 2714 2840
rect -3006 -2880 2714 -2840
rect 3326 2840 9046 2880
rect 3326 -2840 3366 2840
rect 9006 -2840 9046 2840
rect 3326 -2880 9046 -2840
rect -9338 -3240 -3618 -3200
rect -9338 -8920 -9298 -3240
rect -3658 -8920 -3618 -3240
rect -9338 -8960 -3618 -8920
rect -3006 -3240 2714 -3200
rect -3006 -8920 -2966 -3240
rect 2674 -8920 2714 -3240
rect -3006 -8960 2714 -8920
rect 3326 -3240 9046 -3200
rect 3326 -8920 3366 -3240
rect 9006 -8920 9046 -3240
rect 3326 -8960 9046 -8920
<< mimcapcontact >>
rect -9298 3240 -3658 8920
rect -2966 3240 2674 8920
rect 3366 3240 9006 8920
rect -9298 -2840 -3658 2840
rect -2966 -2840 2674 2840
rect 3366 -2840 9006 2840
rect -9298 -8920 -3658 -3240
rect -2966 -8920 2674 -3240
rect 3366 -8920 9006 -3240
<< metal4 >>
rect -6530 8921 -6426 9120
rect -3390 8972 -3286 9120
rect -9299 8920 -3657 8921
rect -9299 3240 -9298 8920
rect -3658 3240 -3657 8920
rect -9299 3239 -3657 3240
rect -6530 2841 -6426 3239
rect -3390 3188 -3370 8972
rect -3306 3188 -3286 8972
rect -198 8921 -94 9120
rect 2942 8972 3046 9120
rect -2967 8920 2675 8921
rect -2967 3240 -2966 8920
rect 2674 3240 2675 8920
rect -2967 3239 2675 3240
rect -3390 2892 -3286 3188
rect -9299 2840 -3657 2841
rect -9299 -2840 -9298 2840
rect -3658 -2840 -3657 2840
rect -9299 -2841 -3657 -2840
rect -6530 -3239 -6426 -2841
rect -3390 -2892 -3370 2892
rect -3306 -2892 -3286 2892
rect -198 2841 -94 3239
rect 2942 3188 2962 8972
rect 3026 3188 3046 8972
rect 6134 8921 6238 9120
rect 9274 8972 9378 9120
rect 3365 8920 9007 8921
rect 3365 3240 3366 8920
rect 9006 3240 9007 8920
rect 3365 3239 9007 3240
rect 2942 2892 3046 3188
rect -2967 2840 2675 2841
rect -2967 -2840 -2966 2840
rect 2674 -2840 2675 2840
rect -2967 -2841 2675 -2840
rect -3390 -3188 -3286 -2892
rect -9299 -3240 -3657 -3239
rect -9299 -8920 -9298 -3240
rect -3658 -8920 -3657 -3240
rect -9299 -8921 -3657 -8920
rect -6530 -9120 -6426 -8921
rect -3390 -8972 -3370 -3188
rect -3306 -8972 -3286 -3188
rect -198 -3239 -94 -2841
rect 2942 -2892 2962 2892
rect 3026 -2892 3046 2892
rect 6134 2841 6238 3239
rect 9274 3188 9294 8972
rect 9358 3188 9378 8972
rect 9274 2892 9378 3188
rect 3365 2840 9007 2841
rect 3365 -2840 3366 2840
rect 9006 -2840 9007 2840
rect 3365 -2841 9007 -2840
rect 2942 -3188 3046 -2892
rect -2967 -3240 2675 -3239
rect -2967 -8920 -2966 -3240
rect 2674 -8920 2675 -3240
rect -2967 -8921 2675 -8920
rect -3390 -9120 -3286 -8972
rect -198 -9120 -94 -8921
rect 2942 -8972 2962 -3188
rect 3026 -8972 3046 -3188
rect 6134 -3239 6238 -2841
rect 9274 -2892 9294 2892
rect 9358 -2892 9378 2892
rect 9274 -3188 9378 -2892
rect 3365 -3240 9007 -3239
rect 3365 -8920 3366 -3240
rect 9006 -8920 9007 -3240
rect 3365 -8921 9007 -8920
rect 2942 -9120 3046 -8972
rect 6134 -9120 6238 -8921
rect 9274 -8972 9294 -3188
rect 9358 -8972 9378 -3188
rect 9274 -9120 9378 -8972
<< properties >>
string FIXED_BBOX 3286 3160 9086 9000
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 28.6 l 28.8 val 1.669k carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
