magic
tech sky130A
magscale 1 2
timestamp 1713418710
<< checkpaint >>
rect 1272 902 4214 1162
rect 1272 690 6374 902
rect 1272 -2778 8220 690
rect 3432 -3038 8220 -2778
rect 5278 -3250 8220 -3038
<< error_s >>
rect 1606 888 1664 894
rect 1606 854 1618 888
rect 1606 848 1664 854
rect 3766 628 3824 634
rect 3766 594 3778 628
rect 3766 588 3824 594
rect 5612 416 5670 422
rect 5612 382 5624 416
rect 5612 376 5670 382
rect 2714 -236 2772 -230
rect 2714 -270 2726 -236
rect 2714 -276 2772 -270
rect 4874 -496 4932 -490
rect 4874 -530 4886 -496
rect 4874 -536 4932 -530
rect 686 -709 739 -708
rect 668 -743 739 -709
rect 669 -744 739 -743
rect 119 -800 200 -777
rect 686 -778 757 -744
rect 1037 -778 1072 -744
rect 147 -828 228 -805
rect 686 -1217 756 -778
rect 1038 -797 1072 -778
rect 868 -846 926 -840
rect 868 -880 880 -846
rect 868 -886 926 -880
rect 868 -1134 926 -1128
rect 868 -1168 880 -1134
rect 868 -1174 926 -1168
rect 686 -1253 739 -1217
rect 1057 -1270 1072 -797
rect 1091 -831 1126 -797
rect 1091 -1270 1125 -831
rect 1237 -899 1295 -893
rect 1237 -933 1249 -899
rect 1237 -939 1295 -933
rect 1237 -1187 1295 -1181
rect 1237 -1221 1249 -1187
rect 1237 -1227 1295 -1221
rect 1091 -1304 1106 -1270
rect 1426 -1323 1441 -797
rect 1460 -1323 1494 -743
rect 1776 -885 1810 -867
rect 1776 -921 1846 -885
rect 1793 -955 1864 -921
rect 1606 -1240 1664 -1234
rect 1606 -1274 1618 -1240
rect 1606 -1280 1664 -1274
rect 1460 -1357 1475 -1323
rect 1793 -1376 1863 -955
rect 1793 -1412 1846 -1376
rect 2534 -1429 2549 -921
rect 2568 -1429 2602 -867
rect 2916 -1257 2954 -936
rect 3197 -1057 3201 -1033
rect 3251 -1221 3255 -1057
rect 3397 -1159 3455 -1153
rect 3397 -1193 3409 -1159
rect 3397 -1199 3455 -1193
rect 2714 -1346 2772 -1340
rect 2714 -1380 2726 -1346
rect 2714 -1386 2772 -1380
rect 2568 -1463 2583 -1429
rect 3215 -1471 3269 -1273
rect 3397 -1447 3455 -1441
rect 3215 -1497 3227 -1471
rect 3217 -1535 3230 -1501
rect 3251 -1569 3264 -1471
rect 3397 -1481 3409 -1447
rect 3397 -1487 3455 -1481
rect 3586 -1583 3601 -1057
rect 3620 -1583 3654 -1003
rect 3936 -1145 3970 -1127
rect 3936 -1181 4006 -1145
rect 3953 -1215 4024 -1181
rect 3766 -1500 3824 -1494
rect 3766 -1534 3778 -1500
rect 3766 -1540 3824 -1534
rect 3620 -1617 3635 -1583
rect 3953 -1636 4023 -1215
rect 3953 -1672 4006 -1636
rect 4694 -1689 4709 -1181
rect 4728 -1689 4762 -1127
rect 5044 -1233 5078 -1215
rect 5044 -1269 5114 -1233
rect 5061 -1303 5132 -1269
rect 4874 -1606 4932 -1600
rect 4874 -1640 4886 -1606
rect 4874 -1646 4932 -1640
rect 4728 -1723 4743 -1689
rect 5061 -1742 5131 -1303
rect 5243 -1371 5301 -1365
rect 5243 -1405 5255 -1371
rect 5243 -1411 5301 -1405
rect 5243 -1659 5301 -1653
rect 5243 -1693 5255 -1659
rect 5243 -1699 5301 -1693
rect 5061 -1778 5114 -1742
rect 5432 -1795 5447 -1269
rect 5466 -1795 5500 -1215
rect 5782 -1357 5816 -1339
rect 5782 -1393 5852 -1357
rect 5799 -1427 5870 -1393
rect 5612 -1712 5670 -1706
rect 5612 -1746 5624 -1712
rect 5612 -1752 5670 -1746
rect 5466 -1829 5481 -1795
rect 5799 -1848 5869 -1427
rect 5799 -1884 5852 -1848
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_sc_hd__inv_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 2954 0 1 -1518
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_MMRDEV  XM1
timestamp 0
transform 1 0 343 0 1 -963
box -396 -290 396 290
use sky130_fd_pr__pfet_01v8_XYUFBL  XM2
timestamp 0
transform 1 0 897 0 1 -1007
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XYUFBL  XM3
timestamp 0
transform 1 0 3426 0 1 -1320
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  XM4
timestamp 0
transform 1 0 3795 0 1 -453
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  XM5
timestamp 0
transform 1 0 4349 0 1 -1435
box -396 -290 396 290
use sky130_fd_pr__nfet_01v8_BBNS5X  XM6
timestamp 0
transform 1 0 4903 0 1 -1068
box -211 -710 211 710
use sky130_fd_pr__pfet_01v8_XYUFBL  XM7
timestamp 0
transform 1 0 5272 0 1 -1532
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  XM8
timestamp 0
transform 1 0 5641 0 1 -665
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  XM9
timestamp 0
transform 1 0 6195 0 1 -1647
box -396 -290 396 290
use sky130_fd_pr__nfet_01v8_BBNS5X  XM10
timestamp 0
transform 1 0 6749 0 1 -1280
box -211 -710 211 710
use sky130_fd_pr__pfet_01v8_XYUFBL  XM11
timestamp 0
transform 1 0 1266 0 1 -1060
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  XM12
timestamp 0
transform 1 0 1635 0 1 -193
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  XM13
timestamp 0
transform 1 0 2189 0 1 -1175
box -396 -290 396 290
use sky130_fd_pr__nfet_01v8_BBNS5X  XM14
timestamp 0
transform 1 0 2743 0 1 -808
box -211 -710 211 710
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vctrl
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vss
port 3 nsew
<< end >>
