magic
tech sky130A
magscale 1 2
timestamp 1713421724
<< error_p >>
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect -29 -178 29 -172
<< pwell >>
rect -216 -300 216 300
<< nmos >>
rect -30 -100 30 100
<< ndiff >>
rect -88 85 -30 100
rect -88 51 -76 85
rect -42 51 -30 85
rect -88 17 -30 51
rect -88 -17 -76 17
rect -42 -17 -30 17
rect -88 -51 -30 -17
rect -88 -85 -76 -51
rect -42 -85 -30 -51
rect -88 -100 -30 -85
rect 30 85 88 100
rect 30 51 42 85
rect 76 51 88 85
rect 30 17 88 51
rect 30 -17 42 17
rect 76 -17 88 17
rect 30 -51 88 -17
rect 30 -85 42 -51
rect 76 -85 88 -51
rect 30 -100 88 -85
<< ndiffc >>
rect -76 51 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -51
rect 42 51 76 85
rect 42 -17 76 17
rect 42 -85 76 -51
<< psubdiff >>
rect -190 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 190 274
rect -190 153 -156 240
rect 156 153 190 240
rect -190 85 -156 119
rect -190 17 -156 51
rect -190 -51 -156 -17
rect -190 -119 -156 -85
rect 156 85 190 119
rect 156 17 190 51
rect 156 -51 190 -17
rect 156 -119 190 -85
rect -190 -240 -156 -153
rect 156 -240 190 -153
rect -190 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 190 -240
<< psubdiffcont >>
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect -190 119 -156 153
rect 156 119 190 153
rect -190 51 -156 85
rect -190 -17 -156 17
rect -190 -85 -156 -51
rect 156 51 190 85
rect 156 -17 190 17
rect 156 -85 190 -51
rect -190 -153 -156 -119
rect 156 -153 190 -119
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -30 100 30 122
rect -30 -122 30 -100
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
<< polycont >>
rect -17 138 17 172
rect -17 -172 17 -138
<< locali >>
rect -190 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 190 274
rect -190 153 -156 240
rect -33 138 -17 172
rect 17 138 33 172
rect 156 153 190 240
rect -190 85 -156 119
rect -190 17 -156 51
rect -190 -51 -156 -17
rect -190 -119 -156 -85
rect -76 85 -42 104
rect -76 17 -42 19
rect -76 -19 -42 -17
rect -76 -104 -42 -85
rect 42 85 76 104
rect 42 17 76 19
rect 42 -19 76 -17
rect 42 -104 76 -85
rect 156 85 190 119
rect 156 17 190 51
rect 156 -51 190 -17
rect 156 -119 190 -85
rect -190 -240 -156 -153
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect 156 -240 190 -153
rect -190 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 190 -240
<< viali >>
rect -17 138 17 172
rect -76 51 -42 53
rect -76 19 -42 51
rect -76 -51 -42 -19
rect -76 -53 -42 -51
rect 42 51 76 53
rect 42 19 76 51
rect 42 -51 76 -19
rect 42 -53 76 -51
rect -17 -172 17 -138
<< metal1 >>
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -82 53 -36 100
rect -82 19 -76 53
rect -42 19 -36 53
rect -82 -19 -36 19
rect -82 -53 -76 -19
rect -42 -53 -36 -19
rect -82 -100 -36 -53
rect 36 53 82 100
rect 36 19 42 53
rect 76 19 82 53
rect 36 -19 82 19
rect 36 -53 42 -19
rect 76 -53 82 -19
rect 36 -100 82 -53
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
<< properties >>
string FIXED_BBOX -173 -257 173 257
<< end >>
