magic
tech sky130A
magscale 1 2
timestamp 1713423503
<< nwell >>
rect 3997 101 4202 399
rect 3982 -458 4309 -304
rect 3982 -602 4310 -458
rect 4000 -626 4310 -602
rect 3988 -1304 4279 -1006
rect 3988 -1306 4078 -1304
<< pwell >>
rect 3962 -178 4088 38
rect 3966 -880 4088 -658
rect 3968 -1594 4086 -1354
<< psubdiff >>
rect 3988 -19 4062 12
rect 3988 -53 4008 -19
rect 4042 -53 4062 -19
rect 3988 -87 4062 -53
rect 3988 -121 4008 -87
rect 4042 -121 4062 -87
rect 3988 -152 4062 -121
rect 3992 -718 4062 -684
rect 3992 -752 4010 -718
rect 4044 -752 4062 -718
rect 3992 -786 4062 -752
rect 3992 -820 4010 -786
rect 4044 -820 4062 -786
rect 3992 -854 4062 -820
rect 3994 -1423 4060 -1380
rect 3994 -1457 4010 -1423
rect 4044 -1457 4060 -1423
rect 3994 -1491 4060 -1457
rect 3994 -1525 4010 -1491
rect 4044 -1525 4060 -1491
rect 3994 -1568 4060 -1525
<< nsubdiff >>
rect 3997 329 4047 363
rect 4081 329 4166 363
rect 4132 301 4166 329
rect 4132 233 4166 267
rect 4132 171 4166 199
rect 3997 137 4047 171
rect 4081 137 4166 171
rect 4104 -378 4154 -344
rect 4188 -378 4273 -344
rect 4239 -406 4273 -378
rect 4239 -474 4273 -440
rect 4239 -536 4273 -508
rect 4104 -570 4154 -536
rect 4188 -570 4273 -536
rect 4074 -1076 4124 -1042
rect 4158 -1076 4243 -1042
rect 4209 -1104 4243 -1076
rect 4209 -1172 4243 -1138
rect 4209 -1234 4243 -1206
rect 4074 -1268 4124 -1234
rect 4158 -1268 4243 -1234
<< psubdiffcont >>
rect 4008 -53 4042 -19
rect 4008 -121 4042 -87
rect 4010 -752 4044 -718
rect 4010 -820 4044 -786
rect 4010 -1457 4044 -1423
rect 4010 -1525 4044 -1491
<< nsubdiffcont >>
rect 4047 329 4081 363
rect 4132 267 4166 301
rect 4132 199 4166 233
rect 4047 137 4081 171
rect 4154 -378 4188 -344
rect 4239 -440 4273 -406
rect 4239 -508 4273 -474
rect 4154 -570 4188 -536
rect 4124 -1076 4158 -1042
rect 4209 -1138 4243 -1104
rect 4209 -1206 4243 -1172
rect 4124 -1268 4158 -1234
<< locali >>
rect 3940 363 4022 380
rect 3940 329 4047 363
rect 4081 329 4166 363
rect 3940 326 4022 329
rect 4132 301 4166 329
rect 4132 233 4166 267
rect 4132 171 4166 199
rect 3798 156 3836 158
rect 3798 122 3800 156
rect 3834 122 3836 156
rect 3997 137 4047 171
rect 4081 137 4166 171
rect 3798 120 3836 122
rect 1708 71 2094 72
rect 1708 37 1709 71
rect 1743 37 2094 71
rect 1708 36 2094 37
rect 2304 59 2348 62
rect 2304 25 2309 59
rect 2343 25 2348 59
rect 2304 22 2348 25
rect 3988 -19 4062 4
rect 3414 -56 3460 -50
rect 3414 -90 3420 -56
rect 3454 -90 3460 -56
rect 3414 -96 3460 -90
rect 3988 -53 4008 -19
rect 4042 -53 4062 -19
rect 3988 -87 4062 -53
rect 3988 -121 4008 -87
rect 4042 -121 4062 -87
rect 3988 -164 4062 -121
rect 1936 -198 2172 -164
rect 3940 -180 4062 -164
rect 3958 -198 4062 -180
rect 1938 -870 1980 -198
rect 3944 -344 4036 -324
rect 3944 -358 4154 -344
rect 4002 -378 4154 -358
rect 4188 -378 4273 -344
rect 4239 -406 4273 -378
rect 4239 -474 4273 -440
rect 4239 -536 4273 -508
rect 3800 -543 3844 -540
rect 3800 -577 3805 -543
rect 3839 -577 3844 -543
rect 4104 -570 4154 -536
rect 4188 -570 4273 -536
rect 3800 -580 3844 -577
rect 2052 -643 2108 -632
rect 2052 -677 2063 -643
rect 2097 -677 2108 -643
rect 2052 -688 2108 -677
rect 2308 -656 2360 -650
rect 2308 -690 2317 -656
rect 2351 -690 2360 -656
rect 2308 -696 2360 -690
rect 3992 -718 4062 -692
rect 3992 -752 4010 -718
rect 4044 -752 4062 -718
rect 3424 -762 3470 -756
rect 3424 -796 3430 -762
rect 3464 -796 3470 -762
rect 3424 -802 3470 -796
rect 3992 -786 4062 -752
rect 3992 -820 4010 -786
rect 4044 -820 4062 -786
rect 3992 -846 4062 -820
rect 1938 -880 2174 -870
rect 1936 -904 2174 -880
rect 3942 -904 4060 -846
rect 1720 -1570 1762 -1568
rect 1936 -1570 1986 -904
rect 3918 -1028 4074 -1024
rect 3950 -1042 4074 -1028
rect 3950 -1058 4124 -1042
rect 3996 -1076 4124 -1058
rect 4158 -1076 4243 -1042
rect 4209 -1104 4243 -1076
rect 4209 -1172 4243 -1138
rect 4209 -1234 4243 -1206
rect 3790 -1246 3836 -1242
rect 3790 -1280 3796 -1246
rect 3830 -1280 3836 -1246
rect 4074 -1268 4124 -1234
rect 4158 -1268 4243 -1234
rect 3790 -1284 3836 -1280
rect 2038 -1344 2102 -1334
rect 2038 -1378 2053 -1344
rect 2087 -1378 2102 -1344
rect 2038 -1388 2102 -1378
rect 2302 -1347 2344 -1344
rect 2302 -1381 2306 -1347
rect 2340 -1381 2344 -1347
rect 2302 -1384 2344 -1381
rect 3994 -1423 4060 -1388
rect 3994 -1457 4010 -1423
rect 4044 -1457 4060 -1423
rect 3410 -1468 3456 -1466
rect 3410 -1502 3416 -1468
rect 3450 -1502 3456 -1468
rect 3410 -1512 3456 -1502
rect 3994 -1491 4060 -1457
rect 3994 -1525 4010 -1491
rect 4044 -1525 4060 -1491
rect 3994 -1566 4060 -1525
rect 1720 -1571 2164 -1570
rect 1720 -1605 1724 -1571
rect 1758 -1605 2164 -1571
rect 3928 -1604 4060 -1566
rect 1720 -1606 2164 -1605
rect 1720 -1608 1762 -1606
rect 1936 -1608 1986 -1606
<< viali >>
rect 3800 122 3834 156
rect 1709 37 1743 71
rect 2309 25 2343 59
rect 3420 -90 3454 -56
rect 3805 -577 3839 -543
rect 2063 -677 2097 -643
rect 2317 -690 2351 -656
rect 3430 -796 3464 -762
rect 3796 -1280 3830 -1246
rect 2053 -1378 2087 -1344
rect 2306 -1381 2340 -1347
rect 3416 -1502 3450 -1468
rect 1724 -1605 1758 -1571
<< metal1 >>
rect 1588 314 2056 410
rect 1588 210 1788 314
rect 1592 71 1792 82
rect 1592 37 1709 71
rect 1743 37 1792 71
rect 1592 -118 1792 37
rect 1868 -298 1908 314
rect 3786 156 3848 164
rect 3786 122 3800 156
rect 3834 122 3848 156
rect 3786 114 3848 122
rect 2290 70 2348 74
rect 3786 70 3846 114
rect 2290 68 3846 70
rect 2290 16 2303 68
rect 2355 16 3846 68
rect 2294 14 3846 16
rect 2348 12 2376 14
rect 4138 -40 4338 38
rect 3396 -46 3478 -42
rect 3396 -98 3411 -46
rect 3463 -98 3478 -46
rect 3396 -102 3478 -98
rect 4138 -92 4175 -40
rect 4227 -92 4338 -40
rect 4138 -162 4338 -92
rect 1868 -304 1912 -298
rect 1868 -384 2126 -304
rect 1868 -1006 1912 -384
rect 3788 -543 3856 -534
rect 3788 -577 3805 -543
rect 3839 -577 3856 -543
rect 3788 -586 3856 -577
rect 2028 -626 2112 -622
rect 2028 -632 2120 -626
rect 2028 -684 2044 -632
rect 2096 -643 2120 -632
rect 2306 -634 2360 -630
rect 3802 -634 3854 -586
rect 2306 -642 3856 -634
rect 2097 -677 2120 -643
rect 2096 -684 2120 -677
rect 2028 -694 2120 -684
rect 2292 -694 2308 -642
rect 2360 -676 3856 -642
rect 2360 -694 3708 -676
rect 2296 -702 3708 -694
rect 3408 -753 3486 -750
rect 3408 -805 3421 -753
rect 3473 -805 3486 -753
rect 3408 -808 3486 -805
rect 4148 -752 4348 -678
rect 4148 -804 4190 -752
rect 4242 -804 4348 -752
rect 4148 -878 4348 -804
rect 1870 -1008 1912 -1006
rect 1870 -1088 2146 -1008
rect 3778 -1246 3848 -1236
rect 3778 -1280 3796 -1246
rect 3830 -1280 3848 -1246
rect 3778 -1290 3848 -1280
rect 2020 -1328 2108 -1326
rect 2020 -1334 2114 -1328
rect 2020 -1386 2038 -1334
rect 2090 -1386 2114 -1334
rect 2290 -1340 2356 -1338
rect 2020 -1394 2114 -1386
rect 2288 -1342 3668 -1340
rect 3790 -1342 3836 -1290
rect 2288 -1347 3838 -1342
rect 2288 -1381 2306 -1347
rect 2340 -1381 3838 -1347
rect 2288 -1390 3838 -1381
rect 2288 -1392 3668 -1390
rect 1590 -1571 1792 -1432
rect 4158 -1452 4358 -1382
rect 3398 -1458 3468 -1452
rect 3388 -1510 3404 -1458
rect 3456 -1510 3472 -1458
rect 4158 -1504 4202 -1452
rect 4254 -1504 4358 -1452
rect 1590 -1605 1724 -1571
rect 1758 -1605 1792 -1571
rect 4158 -1582 4358 -1504
rect 1590 -1634 1792 -1605
<< via1 >>
rect 2303 59 2355 68
rect 2303 25 2309 59
rect 2309 25 2343 59
rect 2343 25 2355 59
rect 2303 16 2355 25
rect 3411 -56 3463 -46
rect 3411 -90 3420 -56
rect 3420 -90 3454 -56
rect 3454 -90 3463 -56
rect 3411 -98 3463 -90
rect 4175 -92 4227 -40
rect 2044 -643 2096 -632
rect 2044 -677 2063 -643
rect 2063 -677 2096 -643
rect 2044 -684 2096 -677
rect 2308 -656 2360 -642
rect 2308 -690 2317 -656
rect 2317 -690 2351 -656
rect 2351 -690 2360 -656
rect 2308 -694 2360 -690
rect 3421 -762 3473 -753
rect 3421 -796 3430 -762
rect 3430 -796 3464 -762
rect 3464 -796 3473 -762
rect 3421 -805 3473 -796
rect 4190 -804 4242 -752
rect 2038 -1344 2090 -1334
rect 2038 -1378 2053 -1344
rect 2053 -1378 2087 -1344
rect 2087 -1378 2090 -1344
rect 2038 -1386 2090 -1378
rect 3404 -1468 3456 -1458
rect 3404 -1502 3416 -1468
rect 3416 -1502 3450 -1468
rect 3450 -1502 3456 -1468
rect 3404 -1510 3456 -1502
rect 4202 -1504 4254 -1452
<< metal2 >>
rect 2300 68 2358 78
rect 2300 16 2303 68
rect 2355 48 2358 68
rect 2355 16 2360 48
rect 2300 -244 2360 16
rect 3406 -44 3468 -32
rect 4174 -40 4228 -24
rect 4174 -44 4175 -40
rect 3406 -46 4175 -44
rect 3406 -98 3411 -46
rect 3463 -92 4175 -46
rect 4227 -92 4228 -40
rect 3463 -98 3468 -92
rect 3406 -112 3468 -98
rect 4174 -108 4228 -92
rect 2040 -294 2360 -244
rect 2040 -612 2102 -294
rect 2038 -632 2102 -612
rect 2038 -684 2044 -632
rect 2096 -684 2102 -632
rect 2038 -704 2102 -684
rect 2302 -642 2366 -632
rect 2302 -694 2308 -642
rect 2360 -694 2366 -642
rect 2302 -704 2366 -694
rect 2306 -948 2364 -704
rect 3418 -752 3476 -740
rect 4188 -750 4244 -730
rect 4090 -752 4244 -750
rect 3418 -753 4190 -752
rect 3418 -805 3421 -753
rect 3473 -804 4190 -753
rect 4242 -804 4244 -752
rect 3473 -805 4244 -804
rect 3418 -808 4244 -805
rect 3418 -818 3476 -808
rect 4188 -826 4244 -808
rect 2044 -988 2364 -948
rect 2044 -1316 2088 -988
rect 2030 -1334 2098 -1316
rect 2030 -1386 2038 -1334
rect 2090 -1386 2098 -1334
rect 2030 -1404 2098 -1386
rect 4196 -1446 4260 -1436
rect 3398 -1452 4262 -1446
rect 3398 -1458 4202 -1452
rect 3398 -1510 3404 -1458
rect 3456 -1504 4202 -1458
rect 4254 -1504 4262 -1452
rect 3456 -1510 4262 -1504
rect 3398 -1520 3462 -1510
rect 4196 -1520 4260 -1510
use sky130_fd_sc_hd__dfxbp_2  x1
timestamp 1713423503
transform 1 0 2032 0 1 -886
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_2  x2
timestamp 1713423503
transform 1 0 2020 0 1 -1588
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_2  x3
timestamp 1713423503
transform 1 0 2028 0 1 -182
box -38 -48 1970 592
<< labels >>
flabel metal1 s 1592 -118 1792 82 0 FreeSans 320 0 0 0 clock
port 1 nsew
flabel metal1 s 4138 -162 4338 38 0 FreeSans 320 0 0 0 out_a
port 2 nsew
flabel metal1 s 4148 -878 4348 -678 0 FreeSans 320 0 0 0 out_b
port 3 nsew
flabel metal1 s 4158 -1582 4358 -1382 0 FreeSans 320 0 0 0 out_c
port 4 nsew
flabel metal1 s 1588 210 1788 410 0 FreeSans 320 0 0 0 vdd
port 5 nsew
flabel metal1 s 1590 -1634 1790 -1434 0 FreeSans 320 0 0 0 vss
port 6 nsew
<< end >>
