magic
tech sky130A
timestamp 1709187259
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
use inverter  x1
timestamp 1709187100
transform 1 0 -259 0 1 -79
box 259 -521 866 29
use inverter  x2
timestamp 1709187100
transform 1 0 348 0 1 -79
box 259 -521 866 29
use inverter  x3
timestamp 1709187100
transform 1 0 955 0 1 -79
box 259 -521 866 29
use inverter31  x31 ~/.xschem/simulations
timestamp 1709187259
transform 1 0 1840 0 1 24
box 69 -764 819 -95
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 inp
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 out
port 3 nsew
<< end >>
