* NGSPICE file created from pfd.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N a_1462_47#
+ a_543_47# a_651_413# a_193_47# a_805_47# a_448_47# a_639_47# a_1283_21# a_761_289#
+ a_1108_47# a_1217_47# a_1659_47# a_1270_413# a_27_47#
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 Q_N a_1659_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.155 ps=1.31 w=1 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR a_1283_21# a_1659_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1522 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 VGND a_1283_21# a_1659_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 VPWR a_1659_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X18 VGND a_1659_47# Q_N VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X20 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X21 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1197 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X26 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10025 ps=0.985 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X29 Q_N a_1659_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.1522 ps=1.335 w=1 l=0.15
X31 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X32 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X33 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X34 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
C0 a_448_47# a_193_47# 0.064178f
C1 Q_N VGND 0.142765f
C2 VPWR Q 0.014118f
C3 RESET_B a_1108_47# 0.236601f
C4 Q_N a_193_47# 9.35e-20
C5 a_1217_47# a_1108_47# 0.007416f
C6 a_761_289# a_639_47# 3.16e-19
C7 VPB a_1659_47# 0.073099f
C8 a_27_47# a_1659_47# 5.63e-20
C9 VGND a_639_47# 0.008634f
C10 a_1283_21# a_543_47# 3.83e-21
C11 VPB a_761_289# 0.099418f
C12 a_1283_21# VPWR 0.156931f
C13 VGND a_1462_47# 0.002121f
C14 a_193_47# a_639_47# 2.28e-19
C15 RESET_B a_1659_47# 0.00263f
C16 a_761_289# a_27_47# 0.07009f
C17 a_448_47# a_543_47# 0.049827f
C18 a_448_47# VPWR 0.068142f
C19 a_1108_47# a_1659_47# 0.00277f
C20 VPB VGND 0.013806f
C21 RESET_B a_761_289# 0.166114f
C22 D a_1283_21# 2.77e-22
C23 a_1217_47# a_761_289# 4.2e-19
C24 VPB a_193_47# 0.170861f
C25 VGND a_27_47# 0.253971f
C26 Q_N VPWR 0.157089f
C27 a_761_289# a_1108_47# 0.051162f
C28 a_193_47# a_27_47# 0.906454f
C29 D a_448_47# 0.155634f
C30 VGND RESET_B 0.28755f
C31 a_1283_21# Q 0.053245f
C32 VGND a_1217_47# 9.68e-19
C33 a_193_47# RESET_B 0.026903f
C34 a_193_47# a_1217_47# 2.36e-20
C35 a_543_47# a_639_47# 0.013793f
C36 VGND a_1108_47# 0.147486f
C37 RESET_B a_1270_413# 2.06e-19
C38 a_193_47# a_1108_47# 0.125324f
C39 a_805_47# RESET_B 0.003155f
C40 Q_N Q 0.0061f
C41 a_1270_413# a_1108_47# 0.006453f
C42 VPB CLK 0.069345f
C43 VPB a_651_413# 0.013543f
C44 VPB a_543_47# 0.095793f
C45 CLK a_27_47# 0.233602f
C46 VPB VPWR 0.250676f
C47 a_651_413# a_27_47# 9.73e-19
C48 a_543_47# a_27_47# 0.115353f
C49 VGND a_1659_47# 0.13852f
C50 VPWR a_27_47# 0.152295f
C51 a_448_47# a_1283_21# 1.11e-21
C52 RESET_B CLK 1.09e-19
C53 RESET_B a_651_413# 0.012196f
C54 a_193_47# a_1659_47# 6.89e-19
C55 RESET_B a_543_47# 0.153272f
C56 Q_N a_1283_21# 0.002658f
C57 VGND a_761_289# 0.073384f
C58 RESET_B VPWR 0.065186f
C59 D VPB 0.137565f
C60 a_193_47# a_761_289# 0.186387f
C61 a_1108_47# a_543_47# 7.99e-20
C62 D a_27_47# 0.132849f
C63 VPWR a_1108_47# 0.171084f
C64 a_761_289# a_1270_413# 2.6e-19
C65 VPB Q 0.002023f
C66 D RESET_B 4.72e-19
C67 a_805_47# a_761_289# 3.69e-19
C68 VGND a_193_47# 0.063057f
C69 a_27_47# Q 3.03e-20
C70 a_1283_21# a_1462_47# 0.007399f
C71 RESET_B Q 8.5e-19
C72 VGND a_805_47# 0.00579f
C73 a_193_47# a_1270_413# 1.46e-19
C74 a_448_47# a_639_47# 4.61e-19
C75 VPWR a_1659_47# 0.205837f
C76 VPB a_1283_21# 0.2414f
C77 a_651_413# a_761_289# 0.097745f
C78 a_761_289# a_543_47# 0.209641f
C79 a_1283_21# a_27_47# 0.043643f
C80 a_761_289# VPWR 0.10497f
C81 VPB a_448_47# 0.014137f
C82 VGND CLK 0.017208f
C83 a_1283_21# RESET_B 0.277236f
C84 VGND a_543_47# 0.122935f
C85 a_448_47# a_27_47# 0.093133f
C86 a_193_47# CLK 7.94e-19
C87 Q_N VPB 0.004225f
C88 VGND VPWR 0.096782f
C89 a_193_47# a_651_413# 0.034619f
C90 a_193_47# a_543_47# 0.229804f
C91 a_1659_47# Q 0.185134f
C92 a_1283_21# a_1108_47# 0.245854f
C93 Q_N a_27_47# 1.53e-20
C94 a_193_47# VPWR 0.395736f
C95 a_448_47# RESET_B 2.45e-19
C96 VPWR a_1270_413# 7.19e-19
C97 a_805_47# a_543_47# 0.001705f
C98 Q_N RESET_B 2.83e-19
C99 D VGND 0.051614f
C100 D a_193_47# 0.217945f
C101 Q_N a_1108_47# 1.34e-19
C102 a_27_47# a_639_47# 0.001881f
C103 VGND Q 0.114874f
C104 a_1283_21# a_1659_47# 0.303605f
C105 a_193_47# Q 1.19e-19
C106 RESET_B a_639_47# 9.54e-19
C107 a_651_413# a_543_47# 0.057222f
C108 CLK VPWR 0.017406f
C109 a_1283_21# a_761_289# 3.17e-21
C110 a_651_413# VPWR 0.12856f
C111 RESET_B a_1462_47# 0.002879f
C112 VPWR a_543_47# 0.100285f
C113 VPB a_27_47# 0.261873f
C114 Q_N a_1659_47# 0.145144f
C115 VPB RESET_B 0.138482f
C116 a_1283_21# VGND 0.2208f
C117 D a_543_47# 7.35e-20
C118 RESET_B a_27_47# 0.296336f
C119 a_1283_21# a_193_47# 0.042424f
C120 D VPWR 0.081188f
C121 a_1217_47# a_27_47# 2.56e-19
C122 VPB a_1108_47# 0.111392f
C123 a_448_47# VGND 0.0661f
C124 a_1108_47# a_27_47# 0.102355f
C125 RESET_B a_1217_47# 6.03e-19
C126 Q_N VNB 0.025191f
C127 Q VNB 0.003804f
C128 VGND VNB 1.24553f
C129 VPWR VNB 1.02447f
C130 RESET_B VNB 0.260034f
C131 D VNB 0.159894f
C132 CLK VNB 0.195254f
C133 VPB VNB 2.19949f
C134 a_1659_47# VNB 0.21348f
C135 a_651_413# VNB 0.004694f
C136 a_448_47# VNB 0.013901f
C137 a_1108_47# VNB 0.127984f
C138 a_1283_21# VNB 0.492394f
C139 a_543_47# VNB 0.157869f
C140 a_761_289# VNB 0.120848f
C141 a_193_47# VNB 0.272482f
C142 a_27_47# VNB 0.495595f
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X a_147_75# a_61_75#
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
C0 B VPWR 0.012524f
C1 VPB A 0.08239f
C2 B a_61_75# 0.142002f
C3 X VPWR 0.194597f
C4 B VGND 0.011526f
C5 B VPB 0.064248f
C6 B A 0.096585f
C7 X a_61_75# 0.149596f
C8 X VGND 0.153129f
C9 X VPB 0.005513f
C10 a_147_75# X 5.82e-19
C11 X A 1.84e-19
C12 VPWR a_61_75# 0.158516f
C13 VPWR VGND 0.07134f
C14 B X 0.002798f
C15 VPWR VPB 0.090199f
C16 a_147_75# VPWR 6.31e-19
C17 VPWR A 0.040281f
C18 a_61_75# VGND 0.125003f
C19 a_61_75# VPB 0.087048f
C20 VPB VGND 0.009503f
C21 a_147_75# a_61_75# 0.006569f
C22 a_147_75# VGND 0.004769f
C23 a_61_75# A 0.085863f
C24 VGND A 0.015556f
C25 VGND VNB 0.390327f
C26 X VNB 0.027496f
C27 B VNB 0.111386f
C28 A VNB 0.177011f
C29 VPWR VNB 0.349659f
C30 VPB VNB 0.604764f
C31 a_61_75# VNB 0.263837f
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
C0 A Y 0.359887f
C1 VGND A 0.081909f
C2 VPWR A 0.098226f
C3 VGND Y 0.262586f
C4 A VPB 0.141975f
C5 VPWR Y 0.361779f
C6 VPB Y 0.015896f
C7 VGND VPWR 0.050092f
C8 VGND VPB 0.006668f
C9 VPWR VPB 0.065385f
C10 VGND VNB 0.326816f
C11 Y VNB 0.084947f
C12 VPWR VNB 0.296394f
C13 A VNB 0.451855f
C14 VPB VNB 0.516168f
.ends

.subckt pfd VSS VDD A QA QB B
Xx1 A VDD x4/Y VSS VSS VDD VDD QA x1/Q_N x1/a_1462_47# x1/a_543_47# x1/a_651_413#
+ x1/a_193_47# x1/a_805_47# x1/a_448_47# x1/a_639_47# x1/a_1283_21# x1/a_761_289#
+ x1/a_1108_47# x1/a_1217_47# x1/a_1659_47# x1/a_1270_413# x1/a_27_47# sky130_fd_sc_hd__dfrbp_2
Xx2 QA QB VSS VSS VDD VDD x4/A x2/a_147_75# x2/a_61_75# sky130_fd_sc_hd__and2_2
Xx3 B VDD x4/Y VSS VSS VDD VDD QB x3/Q_N x3/a_1462_47# x3/a_543_47# x3/a_651_413#
+ x3/a_193_47# x3/a_805_47# x3/a_448_47# x3/a_639_47# x3/a_1283_21# x3/a_761_289#
+ x3/a_1108_47# x3/a_1217_47# x3/a_1659_47# x3/a_1270_413# x3/a_27_47# sky130_fd_sc_hd__dfrbp_2
Xx4 x4/A VSS VSS VDD VDD x4/Y sky130_fd_sc_hd__inv_4
C0 x2/a_147_75# VSS 0.001305f
C1 x3/a_27_47# x4/A 0.002794f
C2 x3/a_761_289# x1/a_543_47# 3.92e-20
C3 x3/a_761_289# x1/a_193_47# 8.32e-21
C4 x3/a_193_47# VSS 0.002869f
C5 x1/a_1659_47# x3/a_1659_47# 0.001065f
C6 x3/a_193_47# x1/a_543_47# 4.23e-19
C7 x3/a_193_47# x1/a_193_47# 2.81e-19
C8 VSS x4/A 0.064922f
C9 x1/a_651_413# x4/Y 0.002005f
C10 x4/Y x3/a_1462_47# 6.94e-20
C11 x1/a_543_47# x4/A 7.24e-19
C12 x4/Y x3/a_1283_21# 0.007804f
C13 x4/A x1/a_193_47# 0.002973f
C14 x1/a_1283_21# VDD 0.013028f
C15 x1/a_27_47# x1/a_1283_21# -1.22e-20
C16 x1/Q_N VDD -0.002396f
C17 x3/a_1283_21# x1/a_1108_47# 2.3e-20
C18 x1/Q_N x1/a_27_47# -4.19e-21
C19 x4/Y x3/a_1270_413# 1.87e-19
C20 x3/a_1283_21# QA 0.002893f
C21 QB x1/a_1283_21# 0.003617f
C22 x4/Y x2/a_61_75# 9.55e-19
C23 x3/a_1283_21# x3/a_27_47# -1.22e-20
C24 x1/Q_N QB 7.23e-19
C25 x4/Y x3/a_543_47# 0.019185f
C26 B x4/Y 0.002946f
C27 x1/a_1108_47# x2/a_61_75# 0.00156f
C28 x4/Y x1/a_448_47# 0.006797f
C29 x1/a_1217_47# VDD 2.11e-20
C30 x4/Y x3/a_651_413# 0.008881f
C31 x3/a_1462_47# VSS 1.7e-19
C32 x3/a_1283_21# VSS 0.005368f
C33 x3/Q_N VDD -0.001965f
C34 x3/a_1283_21# x1/a_193_47# 2.6e-20
C35 x3/a_1108_47# x4/A 4.07e-20
C36 QA x2/a_61_75# -7.04e-19
C37 x4/Y VDD 1.068738f
C38 x3/a_761_289# x4/A 0.002138f
C39 x1/a_27_47# x4/Y 0.021492f
C40 B x3/a_27_47# 0.009415f
C41 B A 0.019541f
C42 x1/a_448_47# QA 2.54e-20
C43 x1/a_1108_47# VDD 0.002912f
C44 x3/a_27_47# x1/a_448_47# 1.92e-21
C45 VSS x3/a_1270_413# 3e-20
C46 QB x3/Q_N 0.076678f
C47 VSS x2/a_61_75# 0.044394f
C48 x3/a_193_47# x4/A 6.35e-19
C49 x3/a_543_47# VSS 0.001259f
C50 B VSS 0.003206f
C51 x4/Y QB 0.050631f
C52 VDD QA 0.252484f
C53 x1/a_1659_47# x3/a_1283_21# 9.92e-21
C54 x3/a_543_47# x1/a_543_47# 0.001216f
C55 x3/a_543_47# x1/a_193_47# 3.36e-21
C56 x3/a_27_47# VDD 0.002308f
C57 x4/Y x1/a_639_47# 0.003447f
C58 VSS x3/a_651_413# 1.73e-19
C59 A VDD 0.276941f
C60 x1/a_27_47# QA 5.73e-19
C61 x1/a_27_47# x3/a_27_47# 7.09e-19
C62 x1/a_27_47# A 0.003469f
C63 x4/Y x3/a_1217_47# 9.15e-20
C64 x4/Y x1/a_761_289# 0.011692f
C65 VSS VDD 1.455216f
C66 x1/a_1270_413# VDD 1.52e-20
C67 QB QA 0.060347f
C68 x1/a_543_47# VDD 0.006114f
C69 x1/a_27_47# VSS 2.8e-19
C70 x1/a_193_47# VDD 0.016797f
C71 x3/a_27_47# QB 6.7e-19
C72 x1/a_27_47# x1/a_543_47# -7.77e-20
C73 x1/a_805_47# VDD 1.49e-19
C74 x1/a_761_289# QA 3.76e-19
C75 x1/a_651_413# x4/A 5.44e-20
C76 VSS QB 0.070345f
C77 x3/a_1108_47# x2/a_61_75# 0.001741f
C78 VSS x1/a_639_47# 1.17e-19
C79 x3/a_1283_21# x4/A 1.74e-19
C80 x3/a_448_47# B 8.04e-20
C81 x1/a_1659_47# VDD 0.003868f
C82 x4/Y x1/a_1283_21# 0.002474f
C83 x1/a_1659_47# x1/a_27_47# -2.46e-20
C84 B x3/a_761_289# 1.38e-19
C85 x3/a_1217_47# VSS 5.01e-20
C86 VSS x1/a_761_289# -0.001714f
C87 x3/a_1659_47# VDD -4.15e-19
C88 x1/Q_N x4/Y 1.8e-19
C89 x4/A x2/a_61_75# 0.0135f
C90 x3/a_1108_47# VDD 5.48e-19
C91 x3/a_193_47# B 0.001165f
C92 x3/a_448_47# VDD 7.49e-20
C93 VDD x1/a_1462_47# 2.14e-20
C94 x3/a_543_47# x4/A 0.001072f
C95 x1/a_27_47# x3/a_1108_47# 2.65e-20
C96 x1/a_1659_47# QB 0.002508f
C97 x3/a_193_47# x1/a_448_47# 2.61e-20
C98 x3/a_761_289# VDD 1.79e-20
C99 x1/a_1283_21# QA 0.025993f
C100 x2/a_147_75# VDD -1.99e-19
C101 x4/A x3/a_651_413# 3.63e-19
C102 QB x3/a_1659_47# 0.096601f
C103 x1/Q_N QA 0.066369f
C104 x3/a_193_47# VDD 0.003037f
C105 x4/Y x1/a_1217_47# 3.35e-19
C106 x3/a_1108_47# QB 0.003568f
C107 x3/a_448_47# QB 2.37e-20
C108 x3/a_193_47# x1/a_27_47# 0.001366f
C109 x4/Y x3/Q_N 5.72e-19
C110 x4/A VDD 0.191959f
C111 VSS x1/a_1283_21# 0.001115f
C112 x3/a_761_289# QB 3.38e-19
C113 x1/a_27_47# x4/A 0.002565f
C114 x1/Q_N VSS 0.00477f
C115 x2/a_147_75# QB 0.002256f
C116 x1/Q_N x1/a_193_47# 1.39e-35
C117 x3/a_193_47# QB 7.35e-19
C118 x4/Y x1/a_1108_47# 0.005587f
C119 x3/a_1283_21# x2/a_61_75# 8.96e-19
C120 x1/a_651_413# x3/a_543_47# 1.24e-21
C121 QB x4/A 0.029153f
C122 x3/a_27_47# x3/Q_N -4.19e-21
C123 x4/Y QA 0.007569f
C124 x1/a_1659_47# x1/a_1283_21# -5.68e-32
C125 x3/a_193_47# x1/a_761_289# 1.78e-20
C126 x4/Y x3/a_27_47# 0.063841f
C127 x4/Y A 2.55e-19
C128 x1/a_1217_47# VSS 5.78e-20
C129 x4/A x1/a_761_289# 0.002468f
C130 VSS x3/Q_N 0.009158f
C131 x3/a_1659_47# x1/a_1283_21# 1.13e-19
C132 x1/a_1108_47# QA 0.002062f
C133 x1/a_651_413# VDD 4.53e-19
C134 x3/a_27_47# x1/a_1108_47# 2.11e-20
C135 x3/a_1283_21# VDD 3.46e-19
C136 x1/Q_N x3/a_1659_47# 2.7e-20
C137 x1/a_27_47# x3/a_1283_21# 4.6e-20
C138 x4/Y VSS 0.55527f
C139 x3/a_1108_47# x1/a_1283_21# 1.76e-20
C140 x4/Y x1/a_543_47# 0.014551f
C141 x4/Y x1/a_193_47# 0.013597f
C142 B x3/a_543_47# 1.13e-19
C143 VSS x1/a_1108_47# 4.55e-19
C144 x3/a_27_47# A 5.05e-19
C145 x4/Y x1/a_805_47# 0.001847f
C146 x1/a_1108_47# x1/a_193_47# 1.42e-32
C147 VDD x3/a_1270_413# 3.44e-21
C148 x3/a_1283_21# QB 0.036568f
C149 VDD x2/a_61_75# 0.015492f
C150 VSS QA 0.079436f
C151 x1/a_1659_47# x3/Q_N 5.94e-20
C152 x3/a_543_47# VDD 0.001555f
C153 x3/a_27_47# VSS 0.001358f
C154 x1/a_543_47# QA 2.62e-19
C155 A VSS 0.003056f
C156 x4/A x1/a_1283_21# 1.59e-19
C157 B VDD 0.037258f
C158 x1/a_193_47# QA 0.001315f
C159 x1/a_27_47# x3/a_543_47# 1.37e-20
C160 x3/a_27_47# x1/a_543_47# 1.11e-21
C161 B x1/a_27_47# 2.72e-20
C162 x3/a_27_47# x1/a_193_47# 5.26e-19
C163 x1/a_448_47# VDD 0.001274f
C164 VDD x3/a_651_413# 4.62e-20
C165 x1/a_1659_47# x4/Y 2.33e-19
C166 QB x3/a_1270_413# 4.92e-20
C167 x4/Y x3/a_1659_47# 0.002286f
C168 QB x2/a_61_75# 0.06191f
C169 VSS x1/a_543_47# -1.78e-19
C170 VSS x1/a_193_47# 2.63e-19
C171 x3/a_543_47# QB 2.49e-19
C172 x3/a_639_47# x4/Y 0.001004f
C173 x1/a_27_47# VDD 0.041518f
C174 x4/Y x3/a_1108_47# 0.015946f
C175 x3/a_448_47# x4/Y 0.006088f
C176 VSS x1/a_805_47# 6.61e-20
C177 x4/Y x1/a_1462_47# 3.98e-19
C178 x4/Y x3/a_805_47# 5.09e-19
C179 x1/a_1659_47# QA 0.084248f
C180 x4/Y x3/a_761_289# 0.028323f
C181 x3/a_1659_47# QA 4.13e-19
C182 x3/a_543_47# x1/a_761_289# 4.26e-20
C183 x3/a_27_47# x3/a_1659_47# -2.46e-20
C184 QB VDD 0.394022f
C185 x1/a_639_47# VDD 3.79e-19
C186 x3/a_193_47# x4/Y 0.078086f
C187 x3/a_1283_21# x1/a_1283_21# 0.001687f
C188 x1/a_1659_47# VSS -2.85e-19
C189 x4/Y x4/A 0.056933f
C190 x3/a_193_47# x1/a_1108_47# 8.83e-21
C191 VSS x3/a_1659_47# 0.006621f
C192 x1/a_1108_47# x4/A 3.75e-19
C193 x1/a_761_289# VDD 0.002021f
C194 x3/a_639_47# VSS 1.05e-19
C195 x1/a_27_47# x1/a_761_289# -2.48e-19
C196 x3/a_1108_47# VSS 0.00166f
C197 VSS x1/a_1462_47# 2.06e-19
C198 VSS x3/a_805_47# 6.63e-20
C199 x3/a_193_47# x3/a_27_47# -1.84e-19
C200 x1/a_1283_21# x2/a_61_75# 8.5e-19
C201 x3/a_1108_47# x1/a_193_47# 2.82e-20
C202 VSS x3/a_761_289# 8.47e-19
C203 x4/A QA 2.26e-20
C204 VDD 0 9.515211f
C205 VSS 0 1.458553f
C206 x4/Y 0 1.310204f
C207 x4/A 0 0.603123f
C208 x3/Q_N 0 0.025191f
C209 QB 0 1.514412f
C210 B 0 0.71044f
C211 x3/a_1659_47# 0 0.21348f
C212 x3/a_651_413# 0 0.004694f
C213 x3/a_448_47# 0 0.013901f
C214 x3/a_1108_47# 0 0.127984f
C215 x3/a_1283_21# 0 0.492394f
C216 x3/a_543_47# 0 0.157869f
C217 x3/a_761_289# 0 0.120848f
C218 x3/a_193_47# 0 0.272482f
C219 x3/a_27_47# 0 0.495595f
C220 QA 0 1.749791f
C221 x2/a_61_75# 0 0.263837f
C222 x1/Q_N 0 0.025191f
C223 A 0 0.706987f
C224 x1/a_1659_47# 0 0.21348f
C225 x1/a_651_413# 0 0.004694f
C226 x1/a_448_47# 0 0.013901f
C227 x1/a_1108_47# 0 0.127984f
C228 x1/a_1283_21# 0 0.492394f
C229 x1/a_543_47# 0 0.157869f
C230 x1/a_761_289# 0 0.120848f
C231 x1/a_193_47# 0 0.272482f
C232 x1/a_27_47# 0 0.495595f
.ends

