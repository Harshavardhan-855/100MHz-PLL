magic
tech sky130A
magscale 1 2
timestamp 1713429292
<< nwell >>
rect 3476 2734 3492 2738
rect 3476 2728 3798 2734
<< locali >>
rect 2164 5434 4264 5444
rect 2164 5378 4274 5434
rect 4080 5326 4274 5378
rect 4080 5276 4084 5326
rect 4002 5214 4084 5276
rect 1358 5114 1504 5162
rect 2358 5124 2504 5172
rect 2846 5112 2992 5160
rect 3266 5114 3412 5162
rect 3686 5120 3832 5168
rect 4000 5150 4084 5214
rect 1070 4810 1122 4818
rect 1070 4776 1079 4810
rect 1113 4776 1122 4810
rect 1070 4768 1122 4776
rect 1358 4512 1410 4922
rect 4126 4498 4272 5148
rect 1002 4312 1150 4316
rect 1000 4272 1150 4312
rect 1000 4268 1148 4272
rect 1360 3662 1412 4072
rect 4116 3938 4272 4498
rect 4116 3928 4268 3938
rect 4126 3652 4268 3928
rect 1006 3420 1154 3464
rect 3112 3267 3882 3274
rect 3112 3233 3834 3267
rect 3868 3233 3882 3267
rect 3112 3226 3882 3233
rect 1358 2812 1410 3222
rect 4116 3082 4268 3652
rect 4120 3080 4268 3082
rect 4120 2810 4266 3080
rect 3742 2712 4266 2810
rect 3434 2664 3476 2668
rect 3434 2630 3438 2664
rect 3472 2630 3476 2664
rect 3434 2626 3476 2630
rect 3742 2628 3778 2712
rect 1004 2572 1152 2616
rect 3110 2440 3234 2480
rect 3432 2382 3480 2570
rect 3900 2382 4078 2422
rect 3430 2296 4078 2382
<< viali >>
rect 4084 5148 4276 5326
rect 1079 4776 1113 4810
rect 3834 3233 3868 3267
rect 3438 2630 3472 2664
rect 3898 2422 4080 2600
<< metal1 >>
rect 4072 5326 4288 5332
rect 1196 5308 1916 5310
rect 1194 5258 1916 5308
rect 2152 5274 3894 5324
rect 1194 5024 1234 5258
rect 2152 5168 2210 5274
rect 1930 5110 2308 5168
rect 4072 5148 4084 5326
rect 4276 5148 4288 5326
rect 4072 5142 4288 5148
rect 4084 5130 4284 5142
rect 3084 5106 3162 5108
rect 3534 5106 3574 5108
rect 3044 5080 3162 5106
rect 1194 4972 1918 5024
rect 922 4826 1122 4910
rect 1236 4826 1286 4972
rect 2298 4970 2364 5020
rect 2984 4970 3050 5020
rect 922 4810 1288 4826
rect 922 4776 1079 4810
rect 1113 4776 1288 4810
rect 922 4768 1288 4776
rect 922 4762 1134 4768
rect 922 4710 1122 4762
rect 1236 4444 1286 4768
rect 1880 4460 1934 4672
rect 3128 4664 3162 5080
rect 3462 5078 3574 5106
rect 3890 5080 4004 5108
rect 3406 4968 3472 5018
rect 3534 4864 3574 5078
rect 3828 4970 3894 5020
rect 3964 4894 4004 5080
rect 3946 4890 4026 4894
rect 3512 4863 3596 4864
rect 3512 4811 3528 4863
rect 3580 4811 3596 4863
rect 3946 4838 3960 4890
rect 4012 4838 4026 4890
rect 3946 4834 4026 4838
rect 3512 4810 3596 4811
rect 1870 4452 1946 4460
rect 1236 4406 1286 4410
rect 1870 4400 1882 4452
rect 1934 4400 1946 4452
rect 1870 4392 1946 4400
rect 2908 4398 2956 4610
rect 4026 4604 4076 4670
rect 1720 4260 1756 4264
rect 1572 4224 1756 4260
rect 1186 3578 1236 4158
rect 1720 4136 1756 4224
rect 1880 4182 1934 4392
rect 2906 4352 4092 4398
rect 2908 4242 2956 4352
rect 3006 4182 3056 4248
rect 1968 4136 2022 4164
rect 1720 4108 2022 4136
rect 1754 4106 2022 4108
rect 1576 3378 1764 3414
rect 1182 2728 1232 3308
rect 1728 3266 1764 3378
rect 1882 3330 1936 3824
rect 3510 3814 3531 3866
rect 3583 3814 3604 3866
rect 2912 3540 2958 3764
rect 4026 3758 4092 4352
rect 4028 3756 4078 3758
rect 4026 3540 4114 3542
rect 2912 3494 4114 3540
rect 2912 3392 2958 3494
rect 3010 3332 3060 3398
rect 1984 3266 2014 3322
rect 3810 3280 3892 3288
rect 1726 3236 2014 3266
rect 3808 3275 3894 3280
rect 3808 3223 3825 3275
rect 3877 3223 3894 3275
rect 3808 3220 3894 3223
rect 3810 3210 3892 3220
rect 3844 3029 3928 3038
rect 1576 2528 1768 2564
rect 1732 2416 1768 2528
rect 1882 2486 1934 2978
rect 3844 2977 3860 3029
rect 3912 2977 3928 3029
rect 3844 2968 3928 2977
rect 2910 2836 2956 2916
rect 4026 2910 4114 3494
rect 4320 3269 4520 3338
rect 4320 3217 4376 3269
rect 4428 3217 4520 3269
rect 4320 3138 4520 3217
rect 2910 2790 3486 2836
rect 2910 2760 2956 2790
rect 2898 2759 2976 2760
rect 2898 2707 2911 2759
rect 2963 2707 2976 2759
rect 2898 2706 2976 2707
rect 2910 2548 2956 2706
rect 3436 2674 3486 2790
rect 3422 2664 3488 2674
rect 3422 2630 3438 2664
rect 3472 2630 3488 2664
rect 3422 2620 3488 2630
rect 3886 2600 4092 2606
rect 1982 2416 2020 2492
rect 3008 2486 3058 2552
rect 3886 2422 3898 2600
rect 4080 2422 4092 2600
rect 3886 2416 4092 2422
rect 1732 2386 2020 2416
rect 3892 2404 4092 2416
<< via1 >>
rect 3528 4811 3580 4863
rect 3960 4838 4012 4890
rect 1882 4400 1934 4452
rect 3531 3814 3583 3866
rect 3825 3267 3877 3275
rect 3825 3233 3834 3267
rect 3834 3233 3868 3267
rect 3868 3233 3877 3267
rect 3825 3223 3877 3233
rect 3860 2977 3912 3029
rect 4376 3217 4428 3269
rect 2911 2707 2963 2759
<< metal2 >>
rect 3956 4902 4016 4904
rect 3916 4890 4016 4902
rect 3522 4863 3592 4878
rect 3522 4811 3528 4863
rect 3580 4811 3592 4863
rect 1880 4462 1936 4470
rect 1880 4452 2330 4462
rect 1880 4400 1882 4452
rect 1934 4400 2330 4452
rect 1880 4392 2330 4400
rect 1880 4382 1936 4392
rect 2258 2768 2330 4392
rect 3522 3876 3592 4811
rect 3916 4838 3960 4890
rect 4012 4838 4016 4890
rect 3916 4824 4016 4838
rect 3520 3866 3594 3876
rect 3520 3814 3531 3866
rect 3583 3814 3594 3866
rect 3520 3804 3594 3814
rect 3916 3470 3982 4824
rect 3700 3448 3982 3470
rect 3700 3400 3980 3448
rect 3700 3050 3760 3400
rect 3820 3276 3882 3298
rect 4368 3276 4436 3288
rect 3820 3275 4436 3276
rect 3820 3223 3825 3275
rect 3877 3269 4436 3275
rect 3877 3223 4376 3269
rect 3820 3217 4376 3223
rect 4428 3217 4436 3269
rect 3820 3206 4436 3217
rect 3820 3200 3882 3206
rect 4368 3198 4436 3206
rect 3700 3029 3982 3050
rect 3700 2977 3860 3029
rect 3912 2977 3982 3029
rect 3700 2972 3982 2977
rect 3852 2970 3982 2972
rect 3854 2958 3918 2970
rect 2908 2768 2966 2770
rect 2258 2759 2970 2768
rect 2258 2707 2911 2759
rect 2963 2707 2970 2759
rect 2258 2698 2970 2707
rect 2908 2696 2966 2698
use sky130_fd_pr__nfet_01v8_MMRDEV  M1
timestamp 1713428059
transform -1 0 1718 0 -1 5140
box -386 -280 386 280
use sky130_fd_pr__pfet_01v8_XYUFBL  M2
timestamp 1713428059
transform 1 0 2331 0 1 5147
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XYUFBL  M3
timestamp 1713428059
transform 1 0 3439 0 1 5145
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  M4
timestamp 1713428059
transform 0 1 2981 -1 0 3789
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  M5
timestamp 1713428059
transform 1 0 1366 0 1 3444
box -386 -280 386 280
use sky130_fd_pr__nfet_01v8_BBNS5X  M6
timestamp 1713428059
transform 0 1 2472 -1 0 3365
box -201 -700 201 700
use sky130_fd_pr__pfet_01v8_XYUFBL  M7
timestamp 1713428059
transform 1 0 3861 0 1 5147
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  M8
timestamp 1713428059
transform 0 1 2981 -1 0 2943
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  M9
timestamp 1713428059
transform -1 0 1364 0 1 2596
box -386 -280 386 280
use sky130_fd_pr__nfet_01v8_BBNS5X  M10
timestamp 1713428059
transform 0 1 2470 1 0 2519
box -201 -700 201 700
use sky130_fd_pr__pfet_01v8_XYUFBL  M11
timestamp 1713428059
transform 1 0 3017 0 1 5147
box -211 -299 211 299
use sky130_fd_pr__pfet_01v8_XGA8MR  M12
timestamp 1713428059
transform 0 1 2979 -1 0 4637
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_MMRDEV  M13
timestamp 1713428059
transform 1 0 1362 0 1 4292
box -386 -280 386 280
use sky130_fd_pr__nfet_01v8_BBNS5X  M14
timestamp 1713428059
transform 0 1 2468 -1 0 4215
box -201 -700 201 700
use sky130_fd_sc_hd__inv_2  x1
timestamp 1713428059
transform 0 1 3216 -1 0 2692
box -38 -48 314 592
<< labels >>
flabel metal1 s 4320 3138 4520 3338 0 FreeSans 320 0 0 0 vss
port 2 nsew
flabel metal1 s 922 4710 1122 4910 0 FreeSans 320 0 0 0 vctrl
port 3 nsew
flabel metal1 s 3892 2404 4092 2604 0 FreeSans 320 0 0 0 out
port 4 nsew
flabel metal1 s 4084 5130 4284 5330 0 FreeSans 320 180 0 0 vdd
port 1 nsew
<< end >>
