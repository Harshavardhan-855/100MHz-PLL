magic
tech sky130A
timestamp 1709124411
<< end >>
