magic
tech sky130A
magscale 1 2
timestamp 1713423889
<< nwell >>
rect 3704 374 3908 384
rect 3672 328 3908 374
rect 3704 44 3908 328
rect 2376 -702 2832 -372
rect 3426 -696 3632 -370
rect 3674 -1434 3858 -1116
<< pwell >>
rect 3668 -174 3920 8
rect 3408 -908 3634 -760
rect 3678 -1726 3860 -1452
<< psubdiff >>
rect 3694 -32 3894 -18
rect 3694 -134 3743 -32
rect 3845 -134 3894 -32
rect 3694 -148 3894 -134
rect 3434 -817 3608 -786
rect 3434 -851 3470 -817
rect 3504 -851 3538 -817
rect 3572 -851 3608 -817
rect 3434 -882 3608 -851
rect 3704 -1504 3834 -1478
rect 3704 -1674 3718 -1504
rect 3820 -1674 3834 -1504
rect 3704 -1700 3834 -1674
<< nsubdiff >>
rect 3708 281 3796 338
rect 3708 247 3737 281
rect 3771 247 3796 281
rect 3708 198 3796 247
rect 3710 192 3796 198
rect 3498 -501 3586 -444
rect 3498 -535 3527 -501
rect 3561 -535 3586 -501
rect 3498 -584 3586 -535
rect 3500 -590 3586 -584
rect 3690 -1209 3778 -1152
rect 3690 -1243 3719 -1209
rect 3753 -1243 3778 -1209
rect 3690 -1292 3778 -1243
rect 3692 -1298 3778 -1292
<< psubdiffcont >>
rect 3743 -134 3845 -32
rect 3470 -851 3504 -817
rect 3538 -851 3572 -817
rect 3718 -1674 3820 -1504
<< nsubdiffcont >>
rect 3737 247 3771 281
rect 3527 -535 3561 -501
rect 3719 -1243 3753 -1209
<< locali >>
rect 3658 312 3772 346
rect 1750 256 1814 312
rect 3737 281 3771 312
rect 3737 196 3771 247
rect 3312 118 3376 122
rect 890 104 1560 106
rect 752 96 1560 104
rect 752 -10 758 96
rect 936 -10 1560 96
rect 3312 84 3327 118
rect 3361 84 3376 118
rect 3312 46 3376 84
rect 3312 12 3327 46
rect 3361 12 3376 46
rect 3312 8 3376 12
rect 752 -16 1560 -10
rect 752 -18 942 -16
rect 3702 -32 3886 -18
rect 3702 -48 3743 -32
rect 3698 -80 3743 -48
rect 3845 -80 3886 -32
rect 3698 -114 3702 -80
rect 3736 -114 3743 -80
rect 3845 -114 3846 -80
rect 3880 -114 3886 -80
rect 3698 -134 3743 -114
rect 3845 -134 3886 -114
rect 3698 -146 3886 -134
rect 3702 -148 3886 -146
rect 3294 -430 3558 -388
rect 3484 -436 3558 -430
rect 3484 -470 3562 -436
rect 3527 -501 3561 -470
rect 3527 -586 3561 -535
rect 4078 -626 4094 -572
rect 1706 -662 1852 -656
rect 1706 -670 1982 -662
rect 1706 -776 1726 -670
rect 1832 -776 1982 -670
rect 2648 -692 2816 -690
rect 3142 -692 3210 -678
rect 2648 -702 3012 -692
rect 2282 -705 3012 -702
rect 2282 -739 2679 -705
rect 2713 -739 2751 -705
rect 2785 -739 3012 -705
rect 2282 -744 3012 -739
rect 3142 -726 3159 -692
rect 3193 -726 3210 -692
rect 3142 -740 3210 -726
rect 3338 -738 4094 -626
rect 2282 -746 2836 -744
rect 2964 -746 3012 -744
rect 2282 -752 2816 -746
rect 4078 -750 4094 -738
rect 4272 -750 4288 -572
rect 2648 -754 2816 -752
rect 1706 -780 1982 -776
rect 3438 -778 3606 -776
rect 1706 -790 1852 -780
rect 3438 -884 3469 -778
rect 3575 -884 3606 -778
rect 3438 -886 3606 -884
rect 1704 -1226 1766 -1168
rect 3548 -1172 3756 -1134
rect 3674 -1178 3754 -1172
rect 3719 -1209 3753 -1178
rect 3719 -1294 3753 -1243
rect 712 -1374 878 -1372
rect 712 -1387 1470 -1374
rect 712 -1493 742 -1387
rect 848 -1493 1470 -1387
rect 712 -1502 1470 -1493
rect 3266 -1377 3324 -1366
rect 3266 -1411 3278 -1377
rect 3312 -1411 3324 -1377
rect 3266 -1449 3324 -1411
rect 3266 -1483 3278 -1449
rect 3312 -1483 3324 -1449
rect 3266 -1494 3324 -1483
rect 712 -1508 878 -1502
rect 3704 -1504 3834 -1486
rect 3704 -1522 3718 -1504
rect 3700 -1524 3718 -1522
rect 3820 -1522 3834 -1504
rect 3820 -1524 3836 -1522
rect 3700 -1702 3715 -1524
rect 3821 -1702 3836 -1524
rect 3700 -1704 3836 -1702
<< viali >>
rect 758 -10 936 96
rect 3327 84 3361 118
rect 3327 12 3361 46
rect 3702 -114 3736 -80
rect 3774 -114 3808 -80
rect 3846 -114 3880 -80
rect 1726 -776 1832 -670
rect 2679 -739 2713 -705
rect 2751 -739 2785 -705
rect 3159 -726 3193 -692
rect 4094 -750 4272 -572
rect 3469 -817 3575 -778
rect 3469 -851 3470 -817
rect 3470 -851 3504 -817
rect 3504 -851 3538 -817
rect 3538 -851 3572 -817
rect 3572 -851 3575 -817
rect 3469 -884 3575 -851
rect 742 -1493 848 -1387
rect 3278 -1411 3312 -1377
rect 3278 -1483 3312 -1449
rect 3715 -1674 3718 -1524
rect 3718 -1674 3820 -1524
rect 3820 -1674 3821 -1524
rect 3715 -1702 3821 -1674
<< metal1 >>
rect 1132 378 1374 608
rect 1132 280 1534 378
rect 696 110 896 154
rect 696 96 954 110
rect 696 -10 758 96
rect 936 -10 954 96
rect 696 -24 954 -10
rect 696 -46 896 -24
rect 1132 -340 1374 280
rect 3306 132 3382 134
rect 4054 132 4254 162
rect 3306 118 4254 132
rect 3306 84 3327 118
rect 3361 84 4254 118
rect 3306 46 4254 84
rect 3306 12 3327 46
rect 3361 12 4254 46
rect 3306 4 4254 12
rect 3306 -4 3382 4
rect 2421 -35 2533 -28
rect 2421 -87 2451 -35
rect 2503 -87 2533 -35
rect 4054 -38 4254 4
rect 2421 -94 2533 -87
rect 3658 -80 3966 -42
rect 3658 -114 3702 -80
rect 3736 -114 3774 -80
rect 3808 -114 3846 -80
rect 3880 -114 3966 -80
rect 3658 -166 3966 -114
rect 3644 -264 3968 -166
rect 1122 -356 1374 -340
rect 1122 -472 1156 -356
rect 1336 -374 1374 -356
rect 1908 -374 2126 -372
rect 1336 -395 2126 -374
rect 1336 -447 1927 -395
rect 1979 -447 1991 -395
rect 2043 -447 2055 -395
rect 2107 -447 2126 -395
rect 1336 -470 2126 -447
rect 2330 -468 2890 -360
rect 1336 -472 1918 -470
rect 1122 -474 1918 -472
rect 1122 -488 1374 -474
rect 1132 -1106 1374 -488
rect 1694 -665 1864 -650
rect 1694 -781 1721 -665
rect 1837 -781 1864 -665
rect 2636 -698 2828 -684
rect 3130 -688 3222 -672
rect 2634 -705 2828 -698
rect 2634 -739 2679 -705
rect 2713 -739 2751 -705
rect 2785 -739 2828 -705
rect 2634 -754 2828 -739
rect 2636 -760 2828 -754
rect 3122 -692 3222 -688
rect 3122 -696 3159 -692
rect 3122 -748 3140 -696
rect 3193 -726 3222 -692
rect 3192 -746 3222 -726
rect 3192 -748 3210 -746
rect 3122 -756 3210 -748
rect 3702 -752 3968 -264
rect 4076 -566 4236 -38
rect 3610 -758 3968 -752
rect 4066 -572 4300 -566
rect 4066 -750 4094 -572
rect 4272 -750 4300 -572
rect 4066 -756 4300 -750
rect 1694 -796 1864 -781
rect 3394 -778 3968 -758
rect 3394 -884 3469 -778
rect 3575 -884 3968 -778
rect 2933 -908 3007 -906
rect 3394 -908 3968 -884
rect 2354 -1016 3968 -908
rect 4138 -948 4338 -920
rect 4108 -964 4338 -948
rect 1132 -1200 1474 -1106
rect 1132 -1208 1374 -1200
rect 3610 -1202 3640 -1102
rect 656 -1366 856 -1330
rect 3260 -1366 3330 -1354
rect 656 -1387 890 -1366
rect 656 -1493 742 -1387
rect 848 -1493 890 -1387
rect 656 -1514 890 -1493
rect 3260 -1372 3666 -1366
rect 3260 -1377 3582 -1372
rect 3260 -1411 3278 -1377
rect 3312 -1411 3582 -1377
rect 3260 -1424 3582 -1411
rect 3634 -1424 3666 -1372
rect 3260 -1436 3666 -1424
rect 3260 -1449 3582 -1436
rect 3260 -1483 3278 -1449
rect 3312 -1483 3582 -1449
rect 3260 -1488 3582 -1483
rect 3634 -1488 3666 -1436
rect 3260 -1492 3666 -1488
rect 3702 -1470 3968 -1016
rect 4028 -981 4338 -964
rect 4028 -1033 4049 -981
rect 4101 -1033 4338 -981
rect 4028 -1045 4338 -1033
rect 4028 -1097 4049 -1045
rect 4101 -1097 4338 -1045
rect 4028 -1114 4338 -1097
rect 4138 -1120 4338 -1114
rect 3702 -1480 3970 -1470
rect 3260 -1506 3330 -1492
rect 3702 -1510 4156 -1480
rect 2502 -1513 2612 -1512
rect 656 -1530 856 -1514
rect 2502 -1565 2531 -1513
rect 2583 -1565 2612 -1513
rect 2502 -1566 2612 -1565
rect 3694 -1524 4156 -1510
rect 3694 -1648 3715 -1524
rect 3626 -1702 3715 -1648
rect 3821 -1702 4156 -1524
rect 3626 -1746 4156 -1702
<< via1 >>
rect 2451 -87 2503 -35
rect 1156 -472 1336 -356
rect 1927 -447 1979 -395
rect 1991 -447 2043 -395
rect 2055 -447 2107 -395
rect 1721 -670 1837 -665
rect 1721 -776 1726 -670
rect 1726 -776 1832 -670
rect 1832 -776 1837 -670
rect 1721 -781 1837 -776
rect 3140 -726 3159 -696
rect 3159 -726 3192 -696
rect 3140 -748 3192 -726
rect 3582 -1424 3634 -1372
rect 3582 -1488 3634 -1436
rect 4049 -1033 4101 -981
rect 4049 -1097 4101 -1045
rect 2531 -1565 2583 -1513
<< metal2 >>
rect 2431 -28 2523 -18
rect 2429 -35 2523 -28
rect 2429 -87 2451 -35
rect 2503 -87 2523 -35
rect 2429 -104 2523 -87
rect 1706 -264 1848 -262
rect 2429 -264 2521 -104
rect 1132 -356 1360 -330
rect 1132 -472 1156 -356
rect 1336 -472 1360 -356
rect 1132 -498 1360 -472
rect 1706 -332 2522 -264
rect 1706 -614 1848 -332
rect 1918 -395 2116 -362
rect 1918 -447 1927 -395
rect 1979 -447 1991 -395
rect 2043 -447 2055 -395
rect 2107 -447 2116 -395
rect 1918 -480 2116 -447
rect 1704 -646 1848 -614
rect 1704 -665 1852 -646
rect 1704 -781 1721 -665
rect 1837 -781 1852 -665
rect 3132 -690 3200 -678
rect 1704 -800 1852 -781
rect 3126 -696 3202 -690
rect 3126 -748 3140 -696
rect 3192 -748 3202 -696
rect 1704 -1034 1840 -800
rect 3126 -988 3202 -748
rect 4038 -974 4112 -954
rect 4006 -981 4112 -974
rect 4006 -988 4049 -981
rect 3126 -1033 4049 -988
rect 4101 -1014 4112 -981
rect 4101 -1033 4134 -1014
rect 1702 -1100 2602 -1034
rect 3126 -1045 4134 -1033
rect 3126 -1088 4049 -1045
rect 3126 -1092 3648 -1088
rect 2514 -1502 2602 -1100
rect 3568 -1358 3648 -1092
rect 4006 -1097 4049 -1088
rect 4101 -1088 4134 -1045
rect 4101 -1097 4112 -1088
rect 4006 -1108 4112 -1097
rect 4038 -1124 4112 -1108
rect 3562 -1372 3654 -1358
rect 3562 -1424 3582 -1372
rect 3634 -1424 3654 -1372
rect 3562 -1436 3654 -1424
rect 3562 -1488 3582 -1436
rect 3634 -1488 3654 -1436
rect 3562 -1502 3654 -1488
rect 2512 -1513 2602 -1502
rect 2512 -1565 2531 -1513
rect 2583 -1565 2602 -1513
rect 2512 -1576 2602 -1565
use sky130_fd_sc_hd__dfrbp_2  x1
timestamp 1713419910
transform 1 0 1478 0 1 -216
box -38 -48 2246 592
use sky130_fd_sc_hd__and2_2  x2
timestamp 1713419910
transform -1 0 3406 0 1 -956
box -38 -48 590 592
use sky130_fd_sc_hd__dfrbp_2  x3
timestamp 1713419910
transform 1 0 1432 0 1 -1698
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_4  x4
timestamp 1713419910
transform -1 0 2372 0 1 -966
box -38 -48 498 592
<< labels >>
flabel metal1 s 1160 394 1360 594 0 FreeSans 320 0 0 0 VDD
port 2 nsew
flabel metal1 s 696 -46 896 154 0 FreeSans 320 0 0 0 A
port 3 nsew
flabel metal1 s 4054 -38 4254 162 0 FreeSans 320 0 0 0 QA
port 4 nsew
flabel metal1 s 656 -1530 856 -1330 0 FreeSans 320 0 0 0 B
port 6 nsew
flabel metal1 s 3922 -1718 4122 -1518 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal1 s 4138 -1120 4338 -920 0 FreeSans 320 0 0 0 QB
port 5 nsew
<< end >>
