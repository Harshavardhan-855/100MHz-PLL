magic
tech sky130A
timestamp 1713418710
<< checkpaint >>
rect -649 -98 1615 -74
rect -649 -122 2600 -98
rect -649 -1654 3585 -122
rect 336 -1678 3585 -1654
rect 1321 -1702 3585 -1678
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
use sky130_fd_sc_hd__dfxbp_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 985 0 1 -1024
box -19 -24 985 296
use sky130_fd_sc_hd__dfxbp_2  x2
timestamp 1712078602
transform 1 0 1970 0 1 -1048
box -19 -24 985 296
use sky130_fd_sc_hd__dfxbp_2  x3
timestamp 1712078602
transform 1 0 0 0 1 -1000
box -19 -24 985 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 b
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 c
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 a
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 vdd
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 vss
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 clk
port 5 nsew
<< end >>
