magic
tech sky130A
magscale 1 2
timestamp 1713421724
<< locali >>
rect 1842 1302 2084 1306
rect 1842 1288 2086 1302
rect 1842 1254 2039 1288
rect 2073 1254 2086 1288
rect 1842 1240 2086 1254
rect 1842 1236 2084 1240
rect 780 900 1042 948
rect 1208 898 1358 944
rect 578 128 726 170
rect 924 128 1072 170
rect 1270 126 1418 168
rect 1962 -56 2156 -40
rect 1962 -90 2107 -56
rect 2141 -90 2156 -56
rect 1962 -104 2156 -90
<< viali >>
rect 2039 1254 2073 1288
rect 2107 -90 2141 -56
<< metal1 >>
rect 280 1222 480 1342
rect 1972 1288 2172 1346
rect 1972 1254 2039 1288
rect 2073 1254 2172 1288
rect 280 1162 786 1222
rect 1036 1168 1418 1224
rect 1652 1219 1748 1232
rect 280 1142 480 1162
rect 1092 1088 1134 1168
rect 1652 1167 1674 1219
rect 1726 1167 1748 1219
rect 1652 1154 1748 1167
rect 1972 1146 2172 1254
rect 284 1011 494 1024
rect 284 959 420 1011
rect 472 959 494 1011
rect 284 946 494 959
rect 284 824 484 946
rect 1412 898 1676 946
rect 1078 786 1150 794
rect 576 782 624 784
rect 576 728 726 782
rect 1078 734 1088 786
rect 1140 734 1150 786
rect 576 356 624 728
rect 1078 726 1150 734
rect 1728 726 1920 768
rect 720 632 784 688
rect 1034 628 1104 684
rect 1352 628 1418 678
rect 1666 628 1736 680
rect 1882 624 1920 726
rect 2008 624 2208 678
rect 1880 566 2208 624
rect 576 302 1498 356
rect 1772 308 1840 360
rect 280 118 480 254
rect 810 226 844 302
rect 1140 260 1212 268
rect 1140 208 1150 260
rect 1202 208 1212 260
rect 1882 258 1920 566
rect 2008 478 2208 566
rect 1848 220 1920 258
rect 1140 200 1212 208
rect 1502 124 1764 168
rect 280 112 490 118
rect 280 60 417 112
rect 469 60 490 112
rect 280 54 490 60
rect 732 -18 1496 36
rect 1758 32 1852 38
rect 1758 -20 1779 32
rect 1831 -20 1852 32
rect 1758 -26 1852 -20
rect 2022 -56 2222 60
rect 2022 -90 2107 -56
rect 2141 -90 2222 -56
rect 2022 -140 2222 -90
<< via1 >>
rect 1674 1167 1726 1219
rect 420 959 472 1011
rect 1088 734 1140 786
rect 1150 208 1202 260
rect 417 60 469 112
rect 1779 -20 1831 32
<< metal2 >>
rect 1662 1232 1738 1242
rect 1658 1219 1738 1232
rect 1658 1167 1674 1219
rect 1726 1167 1738 1219
rect 1658 1144 1738 1167
rect 408 1024 484 1034
rect 1658 1024 1736 1144
rect 408 1011 1736 1024
rect 408 959 420 1011
rect 472 959 1736 1011
rect 408 944 1736 959
rect 408 936 484 944
rect 1088 792 1140 804
rect 1088 786 1204 792
rect 1140 734 1204 786
rect 1088 716 1204 734
rect 1150 260 1204 716
rect 1202 208 1204 260
rect 1150 204 1204 208
rect 1150 190 1202 204
rect 406 124 480 128
rect 406 112 1842 124
rect 406 60 417 112
rect 469 60 1842 112
rect 406 54 1842 60
rect 406 44 480 54
rect 1768 32 1842 54
rect 1768 -20 1779 32
rect 1831 -20 1842 32
rect 1768 -36 1842 -20
use sky130_fd_pr__pfet_01v8_XGAKDL  M1
timestamp 1713421724
transform -1 0 1069 0 1 925
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_PSFW3M  M2
timestamp 1713421724
transform 1 0 1114 0 1 170
box -216 -300 216 300
use sky130_fd_pr__nfet_01v8_PSFW3M  M3
timestamp 1713421724
transform 1 0 768 0 1 170
box -216 -300 216 300
use sky130_fd_pr__pfet_01v8_XGAKDL  M4
timestamp 1713421724
transform 1 0 1385 0 1 925
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_PSFW3M  M5
timestamp 1713421724
transform 1 0 1460 0 1 170
box -216 -300 216 300
use sky130_fd_pr__pfet_01v8_XGAKDL  M6
timestamp 1713421724
transform -1 0 1701 0 1 925
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_PSFW3M  M7
timestamp 1713421724
transform 1 0 1806 0 1 170
box -216 -300 216 300
use sky130_fd_pr__pfet_01v8_XGAKDL  M8
timestamp 1713421724
transform 1 0 753 0 1 925
box -211 -419 211 419
<< labels >>
flabel metal1 s 284 824 484 1024 0 FreeSans 320 0 0 0 qa
port 1 nsew
flabel metal1 s 280 54 480 254 0 FreeSans 320 0 0 0 qb
port 2 nsew
flabel metal1 s 2008 478 2208 678 0 FreeSans 320 0 0 0 cp_out
port 3 nsew
flabel metal1 s 1972 1146 2172 1346 0 FreeSans 320 0 0 0 vdd
port 4 nsew
flabel metal1 s 2022 -140 2222 60 0 FreeSans 320 0 0 0 vss
port 5 nsew
flabel metal1 s 280 1142 480 1342 0 FreeSans 320 0 0 0 cp_bias
port 6 nsew
<< end >>
