magic
tech sky130A
magscale 1 2
timestamp 1713432778
<< pwell >>
rect -307 -2724 307 2724
<< psubdiff >>
rect -271 2654 -175 2688
rect 175 2654 271 2688
rect -271 2592 -237 2654
rect 237 2592 271 2654
rect -271 -2654 -237 -2592
rect 237 -2654 271 -2592
rect -271 -2688 -175 -2654
rect 175 -2688 271 -2654
<< psubdiffcont >>
rect -175 2654 175 2688
rect -271 -2592 -237 2592
rect 237 -2592 271 2592
rect -175 -2688 175 -2654
<< xpolycontact >>
rect -141 2126 141 2558
rect -141 -2558 141 -2126
<< xpolyres >>
rect -141 -2126 141 2126
<< locali >>
rect -271 2654 -175 2688
rect 175 2654 271 2688
rect -271 2592 -237 2654
rect 237 2592 271 2654
rect -271 -2654 -237 -2592
rect 237 -2654 271 -2592
rect -271 -2688 -175 -2654
rect 175 -2688 271 -2654
<< viali >>
rect -125 2143 125 2540
rect -125 -2540 125 -2143
<< metal1 >>
rect -131 2540 131 2552
rect -131 2143 -125 2540
rect 125 2143 131 2540
rect -131 2131 131 2143
rect -131 -2143 131 -2131
rect -131 -2540 -125 -2143
rect 125 -2540 131 -2143
rect -131 -2552 131 -2540
<< properties >>
string FIXED_BBOX -254 -2671 254 2671
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 21.42 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 30.649k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
