** sch_path: /home/vks/pll/xschem/inv.sch
**.subckt inv
x1 out VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_2
x2 net1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__inv_2
x3 net2 VSS VSS VDD VDD out sky130_fd_sc_hd__inv_2
V1 vdd GND vdd
V2 vss GND vss
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.options acct list savecurrents
.temp 25
.param vdd=1.8  vss=0

.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.control
save all
tran 0.1n 0.6u
write inv.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
